* XOR gate implementation using NAND gates

.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include OR.sub
.include XOR.sub
.include FA.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c node_m gnd PULSE(0 1.8 0ns 100ps 100ps 400ns 800ns)
* X1 node_b0 node_m node_b0_in node_x gnd XOR
X1 node_a0 node_b0_in node_m node_c1 node_s0 node_x gnd FA


.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a0) v(node_b0)+2 v(node_b0_in)+4 v(node_m)+6 v(node_s0)+8 v(node_c1)+10
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_cout)+4 v(node_sum)+6
.end
.endc