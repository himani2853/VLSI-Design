* SPICE3 file created from full_adder.ext - technology: scmos
.include TSMC_180nm.txt


.param SUPPLY = 1.8


.global GND

Vdd VDD GND 'SUPPLY'
.option scale=0.09u

V_in_A A gnd PULSE(0 1.8 0ns 100ps 100ps 100ns 200ns)
V_in_B B gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_C C_IN gnd PULSE(0 1.8 0ns 100ps 100ps 250ns 500ns)

M1000 VDD B q1d_2_INPUT_XOR_0/BBAR VDD CMOSP w=4 l=2
+  ad=332 pd=260 as=24 ps=20
M1001 AXORB q1d_2_INPUT_XOR_0/BBAR q1d_2_INPUT_XOR_0/ABAR VDD CMOSP w=4 l=3
+  ad=76 pd=62 as=44 ps=38
M1002 q1d_2_INPUT_XOR_0/BBAR B GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=280 ps=226
M1003 VDD A q1d_2_INPUT_XOR_0/ABAR VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 AXORB B A VDD CMOSP w=4 l=3
+  ad=0 pd=0 as=24 ps=20
M1005 q1d_2_INPUT_XOR_0/ABAR A GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1006 AXORB q1d_2_INPUT_XOR_0/BBAR A Gnd CMOSN w=4 l=3
+  ad=72 pd=60 as=24 ps=20
M1007 AXORB B q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1008 VDD C_IN q1d_2_INPUT_XOR_1/BBAR VDD# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1009 SUM_A_XOR_B_XOR_C q1d_2_INPUT_XOR_1/BBAR q1d_2_INPUT_XOR_1/ABAR VDD CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1010 q1d_2_INPUT_XOR_1/BBAR C_IN GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 VDD AXORB q1d_2_INPUT_XOR_1/ABAR VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 SUM_A_XOR_B_XOR_C C_IN AXORB VDD CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1013 q1d_2_INPUT_XOR_1/ABAR AXORB GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1014 SUM_A_XOR_B_XOR_C q1d_2_INPUT_XOR_1/BBAR AXORB Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1015 SUM_A_XOR_B_XOR_C C_IN q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1016 2_input_OR_0/OUT 2_input_OR_0/A GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1017 2_input_OR_0/a_n7_22# 2_input_OR_0/A VDD VDD CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1018 C_OUT 2_input_OR_0/OUT VDD VDD CMOSP w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1019 C_OUT 2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1020 GND 2_input_OR_0/B 2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 2_input_OR_0/OUT 2_input_OR_0/B 2_input_OR_0/a_n7_22# VDD CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1022 VDD A 2_input_AND_0/OUT VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1023 2_input_AND_0/a_4_n21# B GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1024 2_input_OR_0/B 2_input_AND_0/OUT VDD VDD CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1025 2_input_AND_0/OUT B VDD VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 2_input_OR_0/B 2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1027 2_input_AND_0/OUT A 2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1028 VDD AXORB 2_input_AND_1/OUT VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1029 2_input_AND_1/a_4_n21# C_IN GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1030 2_input_OR_0/A 2_input_AND_1/OUT VDD VDD CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1031 2_input_AND_1/OUT C_IN VDD VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 2_input_OR_0/A 2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1033 2_input_AND_1/OUT AXORB 2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
C0 VDD 2_input_OR_0/A 0.03fF
C1 B A 0.75fF
C2 q1d_2_INPUT_XOR_0/BBAR B 0.03fF
C3 A VDD 0.07fF
C4 B GND 0.18fF
C5 AXORB VDD 0.03fF
C6 2_input_OR_0/A GND 0.44fF
C7 2_input_OR_0/B VDD 0.07fF
C8 2_input_AND_0/OUT A 0.12fF
C9 2_input_OR_0/B 2_input_OR_0/A 0.45fF
C10 VDD# q1d_2_INPUT_XOR_1/BBAR 0.03fF
C11 2_input_AND_0/OUT GND 0.04fF
C12 C_IN SUM_A_XOR_B_XOR_C 0.15fF
C13 B q1d_2_INPUT_XOR_0/ABAR 0.08fF
C14 C_IN q1d_2_INPUT_XOR_1/BBAR 0.03fF
C15 AXORB VDD 0.03fF
C16 AXORB 2_input_AND_1/OUT 0.12fF
C17 2_input_AND_0/OUT 2_input_OR_0/B 0.05fF
C18 AXORB VDD 0.04fF
C19 AXORB A 0.18fF
C20 2_input_AND_1/OUT VDD 0.06fF
C21 AXORB GND 0.33fF
C22 2_input_AND_0/OUT VDD 0.08fF
C23 VDD VDD 0.03fF
C24 VDD VDD 0.03fF
C25 AXORB VDD 0.08fF
C26 VDD A 0.39fF
C27 VDD q1d_2_INPUT_XOR_0/BBAR 0.03fF
C28 2_input_OR_0/OUT C_OUT 0.05fF
C29 AXORB q1d_2_INPUT_XOR_0/ABAR 0.19fF
C30 VDD VDD 0.03fF
C31 2_input_OR_0/B VDD 0.12fF
C32 C_IN q1d_2_INPUT_XOR_1/ABAR 0.51fF
C33 VDD 2_input_OR_0/OUT 0.03fF
C34 AXORB SUM_A_XOR_B_XOR_C 0.18fF
C35 VDD VDD 0.03fF
C36 VDD q1d_2_INPUT_XOR_0/ABAR 0.03fF
C37 VDD 2_input_AND_1/OUT 0.08fF
C38 VDD VDD 0.03fF
C39 A VDD 0.03fF
C40 VDD q1d_2_INPUT_XOR_1/BBAR 0.03fF
C41 2_input_AND_1/OUT GND 0.04fF
C42 VDD q1d_2_INPUT_XOR_0/BBAR 0.09fF
C43 B VDD 0.08fF
C44 SUM_A_XOR_B_XOR_C VDD 0.03fF
C45 A GND 0.11fF
C46 q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C47 C_IN VDD# 0.08fF
C48 C_IN VDD 0.07fF
C49 2_input_OR_0/B GND 0.16fF
C50 AXORB q1d_2_INPUT_XOR_1/ABAR 0.24fF
C51 VDD A 0.08fF
C52 VDD q1d_2_INPUT_XOR_0/ABAR 0.03fF
C53 A q1d_2_INPUT_XOR_0/ABAR 0.11fF
C54 VDD 2_input_OR_0/OUT 0.02fF
C55 q1d_2_INPUT_XOR_0/ABAR GND 0.08fF
C56 B VDD 0.07fF
C57 VDD q1d_2_INPUT_XOR_1/ABAR 0.03fF
C58 VDD 2_input_OR_0/A 0.07fF
C59 SUM_A_XOR_B_XOR_C GND 0.05fF
C60 q1d_2_INPUT_XOR_1/BBAR GND 0.04fF
C61 2_input_OR_0/B VDD 0.03fF
C62 VDD q1d_2_INPUT_XOR_0/ABAR 0.03fF
C63 VDD SUM_A_XOR_B_XOR_C 0.04fF
C64 VDD q1d_2_INPUT_XOR_1/BBAR 0.09fF
C65 2_input_AND_0/OUT VDD 0.03fF
C66 VDD VDD 0.03fF
C67 C_IN AXORB 0.93fF
C68 AXORB VDD 0.07fF
C69 VDD 2_input_OR_0/OUT 0.06fF
C70 AXORB B 0.15fF
C71 VDD VDD# 0.03fF
C72 C_IN VDD 0.12fF
C73 2_input_OR_0/OUT GND 0.15fF
C74 VDD C_OUT 0.03fF
C75 VDD VDD 0.06fF
C76 2_input_OR_0/B 2_input_OR_0/OUT 0.20fF
C77 VDD B 0.14fF
C78 VDD VDD 0.03fF
C79 q1d_2_INPUT_XOR_1/ABAR GND 0.27fF
C80 VDD VDD 0.06fF
C81 C_IN VDD 0.09fF
C82 VDD 2_input_OR_0/A 0.18fF
C83 VDD q1d_2_INPUT_XOR_1/ABAR 0.03fF
C84 q1d_2_INPUT_XOR_1/ABAR VDD 0.03fF
C85 2_input_AND_0/OUT VDD 0.06fF
C86 q1d_2_INPUT_XOR_0/BBAR VDD 0.03fF
C87 VDD 2_input_AND_1/OUT 0.03fF
C88 q1d_2_INPUT_XOR_1/ABAR SUM_A_XOR_B_XOR_C 0.19fF
C89 VDD C_OUT 0.03fF
C90 B VDD 0.09fF
C91 AXORB VDD 0.43fF
C92 C_IN GND 0.17fF
C93 2_input_AND_1/OUT 2_input_OR_0/A 0.05fF
C94 GND C_OUT 0.07fF
C95 2_input_AND_1/OUT Gnd 0.38fF
C96 AXORB Gnd 3.61fF
C97 C_IN Gnd 1.60fF
C98 VDD Gnd 0.56fF
C99 VDD Gnd 0.72fF
C100 2_input_AND_0/OUT Gnd 0.38fF
C101 A Gnd 3.16fF
C102 B Gnd 1.52fF
C103 VDD Gnd 0.56fF
C104 VDD Gnd 0.72fF
C105 GND Gnd 0.66fF
C106 C_OUT Gnd 0.19fF
C107 2_input_OR_0/OUT Gnd 0.41fF
C108 2_input_OR_0/B Gnd 0.52fF
C109 2_input_OR_0/A Gnd 0.78fF
C110 VDD Gnd 0.60fF
C111 VDD Gnd 0.73fF
C112 q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C113 q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C114 SUM_A_XOR_B_XOR_C Gnd 0.24fF
C115 VDD Gnd 0.45fF
C116 VDD# Gnd 0.04fF
C117 VDD Gnd 0.08fF
C118 VDD Gnd 0.45fF
C119 q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C120 q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C121 VDD Gnd 0.45fF
C122 VDD Gnd 0.04fF
C123 VDD Gnd 0.08fF
C124 VDD Gnd 0.45fF
.tran 1n 500n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(A) v(B)+2 v(C_IN)+4 
plot v(SUM_A_XOR_B_XOR_C) v(C_OUT)+2 
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_cout)+4 v(node_sum)+6
.end
.endc