.include TSMC_180nm.txt
* .include NAND.sub
.include NOT.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
X1 node_a node_b node_x gnd NOT
X2 node_b node_c node_x gnd NOT
X3 node_c node_a node_x gnd NOT

* Cload node_a gnd 1f
* Cload node_b gnd 1f
* Cload node_c gnd 1f
* * Add wire connection between node_a and node_out
* R_wire node_a node_out 1m  ; Assuming 1 milli-ohm resistance

.tran 1n 50n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a) v(node_b)+2 v(node_c)+4 v(node_out)+6 
* hardcopy image.ps v(node_a) v(node_out)+2 
.end
.endc
