magic
tech scmos
timestamp 1699691262
<< metal1 >>
rect 53 62 68 66
rect 142 61 158 66
rect 236 61 252 66
rect 52 34 59 38
rect 142 33 148 37
rect 235 33 241 37
rect 325 33 333 37
rect -23 27 -16 31
rect 68 26 74 30
rect 161 26 167 30
rect 252 26 257 30
rect -24 20 -15 24
rect 68 19 76 23
rect 162 19 168 23
rect 253 19 259 23
rect 48 8 51 14
rect 138 8 142 13
rect 230 8 234 13
rect 48 3 69 8
rect 138 3 159 8
rect 230 3 250 8
<< m2contact >>
rect 84 63 89 68
rect -11 -2 -6 6
<< metal2 >>
rect -27 69 329 75
rect 84 68 89 69
rect -11 6 -6 7
rect -26 -2 -11 -1
rect -6 -2 324 -1
rect -26 -8 324 -2
use 2_input_AND  2_input_AND_0
timestamp 1699478438
transform 1 0 -15 0 1 34
box -12 -30 69 33
use 2_input_AND  2_input_AND_1
timestamp 1699478438
transform 1 0 75 0 1 33
box -12 -30 69 33
use 2_input_AND  2_input_AND_2
timestamp 1699478438
transform 1 0 168 0 1 33
box -12 -30 69 33
use 2_input_AND  2_input_AND_3
timestamp 1699478438
transform 1 0 259 0 1 33
box -12 -30 69 33
<< labels >>
rlabel metal1 -21 28 -20 29 1 A0
rlabel metal1 -21 21 -20 22 1 B0
rlabel metal1 54 35 56 36 1 A0_B0
rlabel metal1 70 27 71 28 1 A1
rlabel metal1 71 20 72 21 1 B1
rlabel metal1 146 34 147 35 1 A1_B1
rlabel metal1 163 27 164 28 1 A2
rlabel metal1 164 21 165 22 1 B2
rlabel metal1 238 34 239 35 1 A2_B2
rlabel metal1 253 27 255 28 1 A3
rlabel metal1 254 20 256 21 1 B3
rlabel metal1 330 34 331 35 7 A3_B3
rlabel metal2 105 72 106 73 5 VDD
rlabel metal2 81 -5 82 -4 1 GND
<< end >>
