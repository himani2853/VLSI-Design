magic
tech scmos
timestamp 1698924755
<< nwell >>
rect -12 4 14 23
<< ntransistor >>
rect -1 -11 1 -5
<< ptransistor >>
rect -1 11 1 17
<< ndiffusion >>
rect -2 -11 -1 -5
rect 1 -11 2 -5
<< pdiffusion >>
rect -6 16 -1 17
rect -2 12 -1 16
rect -6 11 -1 12
rect 1 11 2 17
<< ndcontact >>
rect -6 -11 -2 -5
rect 2 -11 7 -5
<< pdcontact >>
rect -6 12 -2 16
rect 2 11 7 17
<< polysilicon >>
rect -1 17 1 20
rect -1 3 1 11
rect -2 -1 1 3
rect -1 -5 1 -1
rect -1 -14 1 -11
<< polycontact >>
rect -6 -1 -2 3
<< metal1 >>
rect -12 23 14 29
rect -6 16 -2 23
rect -6 11 -2 12
rect 2 3 7 11
rect -12 -1 -6 3
rect 2 -1 14 3
rect 2 -5 7 -1
rect -6 -17 -2 -11
rect -11 -23 15 -17
<< labels >>
rlabel metal1 -1 26 5 28 5 vdd
rlabel metal1 -10 0 -8 2 3 in
rlabel metal1 9 0 11 2 7 out
rlabel metal1 -2 -22 4 -20 1 gnd
<< end >>
