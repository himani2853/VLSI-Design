magic
tech scmos
timestamp 1701060155
<< metal1 >>
rect -19 80 769 92
rect 167 69 175 80
rect 61 62 81 68
rect 158 64 186 69
rect 259 65 287 70
rect 356 65 384 70
rect 451 67 479 72
rect 553 66 585 72
rect 659 68 691 74
rect 59 34 66 38
rect 156 35 163 39
rect 257 36 265 40
rect 357 36 363 40
rect 450 37 457 41
rect 554 38 561 42
rect 658 39 666 43
rect 766 42 774 46
rect -13 27 -9 31
rect 83 28 88 32
rect 185 29 189 33
rect 283 29 287 33
rect 377 30 383 34
rect 480 31 485 35
rect 587 32 595 36
rect 691 35 698 39
rect -28 20 -8 24
rect 78 21 87 25
rect 179 22 190 26
rect 280 22 288 26
rect 376 23 381 27
rect 475 24 485 28
rect 581 25 593 29
rect 687 28 697 32
rect -28 1 -23 20
rect 552 15 555 18
rect 122 11 154 12
rect 56 5 88 11
rect 122 7 183 11
rect 250 7 282 13
rect 349 7 381 13
rect 447 8 479 14
rect 552 9 584 15
rect 658 13 690 19
rect 113 6 183 7
rect 117 -14 122 6
rect -23 -26 765 -14
<< m2contact >>
rect 73 20 78 25
rect 173 21 179 26
rect 274 20 280 26
rect 368 21 376 27
rect 468 23 475 28
rect 573 23 581 29
rect 679 26 687 33
rect -28 -4 -23 1
<< metal2 >>
rect -28 -35 -23 -4
rect 73 -35 76 20
rect 173 -35 176 21
rect 274 -35 280 20
rect 368 -35 375 21
rect 468 -35 474 23
rect 573 -35 580 23
rect 679 -35 687 26
rect -28 -38 687 -35
use 2_input_AND  2_input_AND_0
timestamp 1699478438
transform 1 0 -7 0 1 34
box -12 -30 69 33
use 2_input_AND  2_input_AND_1
timestamp 1699478438
transform 1 0 90 0 1 35
box -12 -30 69 33
use 2_input_AND  2_input_AND_2
timestamp 1699478438
transform 1 0 191 0 1 36
box -12 -30 69 33
use 2_input_AND  2_input_AND_3
timestamp 1699478438
transform 1 0 290 0 1 36
box -12 -30 69 33
use 2_input_AND  2_input_AND_4
timestamp 1699478438
transform 1 0 384 0 1 37
box -12 -30 69 33
use 2_input_AND  2_input_AND_5
timestamp 1699478438
transform 1 0 487 0 1 38
box -12 -30 69 33
use 2_input_AND  2_input_AND_6
timestamp 1699478438
transform 1 0 593 0 1 39
box -12 -30 69 33
use 2_input_AND  2_input_AND_7
timestamp 1699478438
transform 1 0 699 0 1 42
box -12 -30 69 33
<< labels >>
rlabel metal1 -11 28 -10 29 1 A0
rlabel metal1 695 36 696 37 1 B3
rlabel metal1 588 32 589 34 1 B2
rlabel metal1 481 31 484 32 1 B1
rlabel metal1 379 31 380 32 1 B0
rlabel metal1 284 30 285 31 1 A3
rlabel metal1 187 30 188 31 1 A2
rlabel metal1 84 29 86 30 1 A1
rlabel metal1 64 35 64 36 1 A0_FINAL
rlabel metal1 161 36 162 37 1 A1_FINAL
rlabel metal1 261 37 262 38 1 A2_FINAL
rlabel metal1 360 37 361 38 1 A3_FINAL
rlabel metal1 454 38 455 39 1 B0_FINAL
rlabel metal1 559 40 559 41 1 B1_FINAL
rlabel metal1 658 39 666 43 1 B2_FINAL
rlabel metal1 766 42 774 46 7 B3_FINAL
rlabel metal1 569 -22 572 -21 1 GND
rlabel metal1 559 85 562 86 1 VDD
rlabel metal1 -26 11 -25 12 3 enable
<< end >>
