.include TSMC_180nm.txt
.include 4_input_NOR.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}

.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}


.param wp1 = wn1
.param wp2 = wn1

.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}


.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_b node_b gnd PULSE(0 1.8 0ns 100ps 100ps 160ns 320ns)
V_in_c node_c gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_d node_d gnd PULSE(0 1.8 0ns 100ps 100ps 160ns 320ns)

X1 node_a node_b node_c node_d node_out node_x gnd 4_input_NOR

C1 node_out gnd 100f


.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a) v(node_b)+2 v(node_c)+4 v(node_d)+6 v(node_out)+8
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc