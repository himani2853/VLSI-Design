magic
tech scmos
timestamp 1700304769
<< metal1 >>
rect 1333 181 1659 182
rect 1333 180 1765 181
rect 431 179 1765 180
rect -24 177 1765 179
rect -25 172 1765 177
rect -25 170 1358 172
rect -25 169 455 170
rect -25 154 -15 169
rect -25 150 1 154
rect 61 153 91 169
rect -25 139 -5 150
rect 61 145 62 153
rect -25 137 1 139
rect 191 113 199 169
rect 492 151 515 170
rect 514 144 515 151
rect 902 148 926 170
rect 1037 141 1046 170
rect 1309 156 1327 170
rect 1642 125 1659 172
rect 286 97 295 98
rect -49 87 6 94
rect 278 90 295 97
rect -48 -1 -30 87
rect -25 86 6 87
rect -16 8 11 11
rect -16 0 5 8
rect 155 7 167 15
rect -49 -105 -29 -1
rect -16 -7 11 0
rect -16 -76 -5 -7
rect 157 -10 163 7
rect 206 -16 214 58
rect 190 -27 214 -16
rect 286 -50 295 90
rect 399 94 424 95
rect 399 86 433 94
rect 707 90 720 97
rect 1128 94 1142 96
rect 399 85 424 86
rect 399 45 420 85
rect 399 37 421 45
rect 400 -4 421 37
rect 590 12 595 13
rect 583 7 595 12
rect 400 -16 402 -4
rect 590 -16 595 7
rect 712 -31 720 90
rect 796 85 853 93
rect 1128 89 1149 94
rect 796 84 847 85
rect 796 -7 810 84
rect 1013 11 1020 13
rect 1005 6 1020 11
rect 1013 -10 1020 6
rect 1038 -8 1046 58
rect 1139 -11 1149 89
rect 1233 92 1251 100
rect 1525 96 1526 103
rect 1527 96 1559 103
rect 1570 96 1595 103
rect 1233 32 1250 92
rect 1591 88 1595 96
rect 1697 93 1714 98
rect 1591 84 1611 88
rect 1526 78 1621 81
rect 1527 38 1533 78
rect 1545 72 1628 75
rect 1526 37 1534 38
rect 1404 16 1416 19
rect 1404 11 1420 16
rect 1410 1 1420 11
rect 1441 2 1447 24
rect 1526 21 1535 37
rect 1545 36 1553 72
rect 1571 65 1638 68
rect 1139 -16 1166 -11
rect 1140 -20 1166 -16
rect 1526 -11 1534 21
rect 1180 -20 1534 -11
rect 1545 20 1554 36
rect 1571 35 1579 65
rect 1753 58 1765 172
rect 1571 33 1581 35
rect 1572 24 1581 33
rect 711 -40 734 -31
rect 768 -31 1289 -30
rect 1545 -31 1553 20
rect 751 -39 1553 -31
rect 751 -40 949 -39
rect 1285 -40 1427 -39
rect 1545 -40 1553 -39
rect 1571 19 1581 24
rect 1571 -49 1579 19
rect 1517 -50 1580 -49
rect 286 -59 1580 -50
rect 1617 -60 1628 50
rect 1752 9 1767 58
rect 1934 8 1948 9
rect 1768 -15 1949 8
rect 1615 -75 1628 -60
rect 1483 -76 1628 -75
rect -16 -91 75 -76
rect 103 -91 444 -76
rect -16 -93 444 -91
rect 476 -92 887 -76
rect 898 -91 1289 -76
rect 1324 -84 1628 -76
rect 1324 -91 1747 -84
rect 898 -92 1747 -91
rect 476 -93 821 -92
rect -16 -94 821 -93
rect -47 -147 -30 -105
rect -47 -153 4 -147
rect 24 -153 61 -147
rect 117 -169 126 -94
rect 135 -116 140 -94
rect 183 -130 211 -125
rect 157 -139 161 -135
rect 154 -144 161 -139
rect 146 -170 150 -153
rect 154 -166 158 -144
rect 162 -167 166 -156
rect 178 -160 179 -157
rect 178 -167 182 -160
rect 203 -164 211 -130
rect 567 -124 576 -94
rect 284 -155 285 -148
rect 284 -164 300 -155
rect 177 -617 181 -265
rect 285 -322 299 -164
rect 324 -270 349 -126
rect 552 -152 574 -142
rect 590 -145 595 -141
rect 615 -144 636 -137
rect 992 -123 1000 -92
rect 1398 -93 1747 -92
rect 1421 -112 1489 -104
rect 577 -151 596 -145
rect 552 -190 562 -152
rect 577 -211 581 -151
rect 584 -201 587 -160
rect 590 -191 594 -176
rect 631 -187 636 -144
rect 570 -219 574 -212
rect 733 -240 752 -138
rect 732 -266 752 -240
rect 359 -288 451 -275
rect 324 -290 451 -288
rect 285 -338 382 -322
rect 355 -356 380 -338
rect 356 -375 380 -356
rect 355 -477 380 -375
rect 424 -418 450 -290
rect 598 -358 606 -281
rect 598 -387 606 -386
rect 424 -419 563 -418
rect 732 -419 750 -266
rect 775 -324 785 -162
rect 989 -180 996 -135
rect 1014 -147 1018 -141
rect 1039 -142 1059 -136
rect 1010 -152 1018 -147
rect 1010 -195 1013 -152
rect 1017 -185 1021 -169
rect 1052 -177 1059 -142
rect 1445 -148 1450 -147
rect 1387 -177 1396 -149
rect 1412 -154 1416 -151
rect 1435 -152 1450 -148
rect 1404 -186 1408 -171
rect 1411 -184 1416 -154
rect 1445 -177 1450 -152
rect 1003 -204 1006 -197
rect 1181 -249 1182 -231
rect 1024 -302 1028 -257
rect 1168 -324 1182 -249
rect 775 -346 1182 -324
rect 424 -447 752 -419
rect 424 -449 563 -447
rect 424 -451 450 -449
rect 868 -477 892 -346
rect 1418 -398 1422 -252
rect 1480 -306 1489 -112
rect 1678 -369 1690 -134
rect 1418 -403 1573 -398
rect 1373 -414 1579 -407
rect 1695 -411 1721 -403
rect 1373 -427 1389 -414
rect 1732 -419 1747 -93
rect 1934 -390 1948 -15
rect 1417 -425 1578 -419
rect 1417 -461 1434 -425
rect 1732 -429 1748 -419
rect 1472 -436 1583 -430
rect 355 -506 897 -477
rect 1472 -501 1487 -436
rect 1679 -438 1748 -429
rect 1471 -503 1487 -501
rect 1471 -552 1486 -503
rect 1519 -572 1529 -566
rect 1233 -611 1234 -602
rect 1233 -617 1256 -611
rect 177 -626 1256 -617
rect 1519 -612 1520 -572
rect 177 -627 1246 -626
rect 1419 -731 1424 -687
rect 1441 -713 1445 -693
rect 1519 -695 1529 -612
rect 1733 -695 1748 -438
rect 1934 -549 1950 -390
rect 1936 -657 1950 -549
rect 1519 -707 1520 -695
rect 1731 -730 1748 -695
rect 1831 -730 1862 -728
rect 1723 -731 1862 -730
rect 55 -750 62 -741
rect 78 -742 82 -738
rect 1419 -743 1862 -731
rect 55 -755 909 -750
rect 55 -756 912 -755
rect 57 -833 63 -756
rect 86 -831 90 -774
rect 94 -830 98 -772
rect 102 -786 139 -779
rect 102 -831 106 -786
rect 110 -804 412 -797
rect 110 -830 114 -804
rect 118 -830 122 -817
rect 449 -824 456 -756
rect 902 -775 912 -756
rect 927 -765 931 -751
rect 1424 -765 1440 -743
rect 922 -768 932 -765
rect 1422 -775 1442 -765
rect 535 -788 555 -780
rect 449 -827 474 -824
rect 142 -856 178 -849
rect 468 -850 474 -827
rect 456 -872 473 -865
rect 457 -907 462 -872
rect 489 -877 495 -870
rect 479 -882 495 -877
rect 535 -885 540 -788
rect 902 -785 1442 -775
rect 902 -787 1440 -785
rect 482 -889 542 -885
rect 474 -913 478 -912
rect 116 -928 121 -923
rect 116 -937 122 -928
rect 474 -935 478 -918
rect 482 -926 485 -889
rect 545 -892 551 -820
rect 902 -828 906 -787
rect 923 -842 927 -806
rect 930 -818 1059 -812
rect 930 -833 934 -818
rect 1306 -837 1314 -787
rect 915 -850 919 -843
rect 1306 -845 1426 -837
rect 992 -858 1006 -856
rect 992 -861 995 -858
rect 966 -866 995 -861
rect 1005 -866 1006 -858
rect 488 -895 551 -892
rect 488 -916 491 -895
rect 937 -914 941 -903
rect 116 -1000 121 -937
rect 538 -976 753 -975
rect 992 -976 1006 -866
rect 1419 -923 1425 -845
rect 1474 -852 1486 -781
rect 1540 -790 1727 -773
rect 1435 -863 1486 -852
rect 1435 -931 1439 -863
rect 1708 -870 1727 -790
rect 1442 -875 1727 -870
rect 1442 -877 1726 -875
rect 1442 -930 1446 -877
rect 1831 -890 1862 -743
rect 1477 -924 1483 -892
rect 115 -1056 121 -1000
rect 503 -993 508 -990
rect 538 -993 1006 -976
rect 503 -1004 512 -993
rect 1449 -1001 1453 -999
rect 115 -1185 120 -1056
rect 504 -1120 512 -1004
rect 964 -1120 970 -1119
rect 504 -1127 971 -1120
rect 115 -1198 958 -1185
rect 950 -1205 957 -1198
rect 950 -1212 958 -1205
rect 953 -1338 958 -1212
rect 964 -1341 970 -1127
rect 975 -1340 980 -1033
rect 1448 -1079 1453 -1001
rect 985 -1085 1234 -1084
rect 1448 -1085 1452 -1079
rect 985 -1095 1452 -1085
rect 985 -1203 991 -1095
rect 1827 -1108 1865 -890
rect 1356 -1125 1865 -1108
rect 985 -1223 992 -1203
rect 1357 -1223 1378 -1125
rect 1827 -1126 1865 -1125
rect 986 -1341 992 -1223
rect 1356 -1258 1378 -1223
rect 1356 -1352 1377 -1258
rect 1356 -1370 1378 -1352
rect 910 -1450 922 -1405
rect 909 -1479 922 -1450
rect 978 -1474 986 -1462
rect 909 -1484 923 -1479
rect 1357 -1484 1378 -1370
rect 909 -1498 1378 -1484
rect 1357 -1499 1378 -1498
<< m2contact >>
rect -5 139 2 150
rect 62 142 93 153
rect 492 144 514 151
rect 902 142 926 148
rect 1309 150 1327 156
rect 1037 133 1046 141
rect 191 103 199 113
rect 206 58 215 69
rect 5 0 14 8
rect 157 -18 163 -10
rect 180 -27 190 -15
rect 402 -18 423 -4
rect 590 -22 595 -16
rect 1038 58 1046 68
rect 795 -15 811 -7
rect 1013 -16 1020 -10
rect 1038 -17 1046 -8
rect 1559 96 1570 103
rect 1231 21 1250 32
rect 1441 24 1448 44
rect 1410 -6 1420 1
rect 1436 -5 1447 2
rect 1166 -22 1180 -8
rect 734 -40 751 -29
rect 1752 -15 1768 9
rect 75 -91 103 -76
rect 444 -93 476 -76
rect 887 -92 898 -76
rect 1289 -91 1324 -76
rect 4 -159 24 -146
rect 61 -153 77 -146
rect 156 -114 162 -106
rect 181 -114 192 -108
rect 144 -153 150 -148
rect 161 -156 166 -150
rect 179 -160 185 -155
rect 170 -168 175 -162
rect 324 -126 350 -114
rect 590 -122 595 -116
rect 285 -155 305 -145
rect 731 -138 755 -121
rect 1411 -112 1421 -104
rect 1013 -120 1020 -114
rect 1039 -121 1047 -116
rect 1390 -135 1396 -126
rect 1411 -128 1418 -121
rect 1436 -130 1447 -123
rect 569 -212 574 -207
rect 584 -160 589 -155
rect 590 -176 597 -170
rect 772 -162 786 -152
rect 316 -288 359 -270
rect 598 -386 610 -358
rect 1002 -197 1007 -192
rect 1017 -169 1022 -163
rect 1402 -171 1408 -166
rect 1168 -249 1181 -227
rect 1021 -314 1031 -302
rect 1678 -134 1692 -112
rect 1480 -326 1490 -306
rect 1373 -443 1389 -427
rect 1417 -484 1435 -461
rect 1469 -589 1488 -552
rect 1234 -611 1261 -596
rect 1520 -612 1534 -572
rect 1441 -676 1446 -670
rect 1465 -682 1480 -664
rect 77 -721 83 -710
rect 103 -722 112 -715
rect 927 -735 935 -726
rect 951 -737 958 -729
rect 1920 -684 1957 -657
rect 1520 -707 1529 -695
rect 1441 -718 1447 -713
rect 78 -747 83 -742
rect 85 -774 90 -769
rect 94 -772 104 -765
rect 139 -787 158 -778
rect 412 -804 428 -796
rect 118 -817 127 -811
rect 915 -769 922 -764
rect 178 -857 191 -849
rect 490 -853 496 -842
rect 514 -850 521 -842
rect 474 -882 479 -877
rect 555 -789 564 -779
rect 1473 -781 1486 -765
rect 545 -820 557 -805
rect 474 -918 479 -913
rect 923 -806 932 -795
rect 915 -843 920 -838
rect 1059 -818 1089 -810
rect 995 -866 1005 -858
rect 494 -907 499 -902
rect 937 -921 945 -914
rect 1520 -790 1540 -773
rect 1477 -892 1486 -884
rect 974 -1033 985 -1005
rect 1020 -1440 1041 -1414
<< metal2 >>
rect 225 155 466 162
rect 654 155 894 162
rect 2 139 29 150
rect 447 140 466 155
rect 879 139 893 155
rect 1075 154 1237 161
rect 1230 153 1237 154
rect 1230 146 1289 153
rect 199 103 216 111
rect 206 69 216 103
rect 215 58 216 69
rect 1038 68 1045 133
rect 1441 44 1447 169
rect 1474 161 1475 168
rect 1560 92 1568 96
rect 1510 85 1568 92
rect 1211 21 1231 30
rect 1474 25 1483 32
rect 1211 20 1249 21
rect 14 0 32 8
rect 1254 7 1281 13
rect 1228 6 1281 7
rect 75 -76 103 6
rect 224 0 286 6
rect 295 0 474 6
rect 652 0 877 6
rect 157 -51 162 -18
rect 400 -18 402 -5
rect 157 -106 162 -63
rect 181 -108 189 -27
rect 263 -124 324 -114
rect 263 -138 268 -124
rect 162 -143 268 -138
rect 2 -159 4 -146
rect 24 -159 25 -146
rect 77 -153 144 -148
rect 162 -150 166 -143
rect 170 -151 285 -147
rect 2 -262 25 -159
rect 170 -162 174 -151
rect 400 -153 423 -18
rect 444 -76 474 0
rect 797 -7 810 -6
rect 590 -16 595 -9
rect 590 -98 595 -22
rect 590 -116 595 -110
rect 734 -121 749 -40
rect 797 -145 810 -15
rect 887 -76 898 4
rect 1076 -2 1259 6
rect 1013 -99 1020 -16
rect 985 -105 1020 -99
rect 1013 -114 1020 -105
rect 1038 -116 1046 -17
rect 1180 -22 1181 -9
rect 1038 -121 1039 -116
rect 929 -145 937 -144
rect 185 -160 241 -156
rect 233 -189 241 -160
rect 234 -234 241 -189
rect 401 -198 423 -153
rect 589 -160 648 -155
rect 665 -160 772 -155
rect 797 -157 937 -145
rect 597 -176 704 -170
rect 400 -206 423 -198
rect 400 -211 479 -206
rect 405 -212 479 -211
rect 502 -207 541 -206
rect 502 -212 569 -207
rect 0 -336 26 -262
rect 233 -287 241 -234
rect 233 -290 243 -287
rect -1 -366 26 -336
rect -1 -471 25 -366
rect 234 -405 243 -290
rect 319 -356 357 -288
rect 274 -358 357 -356
rect 263 -371 357 -358
rect 263 -375 356 -371
rect -1 -477 27 -471
rect 1 -578 27 -477
rect 233 -525 245 -405
rect 263 -430 293 -375
rect 679 -367 704 -176
rect 929 -193 937 -157
rect 1089 -162 1103 -159
rect 1017 -163 1103 -162
rect 1022 -169 1103 -163
rect 929 -197 1002 -193
rect 1089 -275 1103 -169
rect 1166 -227 1181 -22
rect 1289 -76 1325 14
rect 1324 -91 1325 -76
rect 1390 -126 1396 12
rect 1411 -104 1419 -6
rect 1411 -121 1419 -112
rect 1418 -128 1419 -121
rect 1436 -123 1447 -5
rect 1510 -23 1523 85
rect 1560 84 1568 85
rect 1379 -171 1402 -166
rect 1166 -245 1168 -227
rect 1509 -203 1523 -23
rect 1678 -13 1752 4
rect 1678 -112 1690 -13
rect 1211 -275 1229 -273
rect 1509 -275 1521 -203
rect 1089 -285 1119 -275
rect 1136 -285 1521 -275
rect 1024 -349 1028 -314
rect 1211 -366 1229 -285
rect 1480 -306 1489 -304
rect 789 -367 1232 -366
rect 598 -447 606 -386
rect 679 -388 1232 -367
rect 679 -389 1122 -388
rect 954 -524 976 -389
rect 1038 -443 1373 -429
rect 1038 -444 1387 -443
rect 1363 -463 1417 -462
rect 1087 -471 1417 -463
rect 303 -525 976 -524
rect 233 -537 976 -525
rect 1085 -483 1417 -471
rect 233 -552 974 -537
rect 233 -553 913 -552
rect 0 -583 84 -578
rect 1085 -582 1104 -483
rect 1363 -484 1417 -483
rect 1480 -466 1489 -326
rect 1519 -466 1529 -465
rect 1480 -474 1529 -466
rect 1236 -573 1469 -564
rect 591 -583 1104 -582
rect 1 -584 27 -583
rect 78 -639 83 -583
rect 615 -598 1104 -583
rect 1235 -587 1469 -573
rect 1235 -596 1254 -587
rect 1519 -572 1529 -474
rect 1519 -606 1520 -572
rect 77 -668 83 -639
rect 513 -646 531 -644
rect 1309 -645 1445 -644
rect 447 -647 993 -646
rect 99 -659 993 -647
rect 1327 -654 1445 -645
rect 99 -666 212 -659
rect 78 -710 83 -668
rect 103 -715 112 -666
rect 227 -665 993 -659
rect 227 -666 621 -665
rect 83 -747 90 -744
rect 86 -769 90 -747
rect 130 -765 137 -705
rect 104 -772 137 -765
rect 139 -778 301 -777
rect 158 -787 260 -778
rect 299 -787 301 -778
rect 490 -790 496 -788
rect 127 -816 350 -811
rect 191 -857 210 -850
rect 413 -1014 425 -804
rect 513 -798 531 -666
rect 555 -779 561 -688
rect 969 -702 993 -665
rect 1441 -670 1445 -654
rect 1632 -661 1660 -660
rect 1919 -661 1920 -658
rect 1465 -664 1920 -661
rect 1480 -682 1920 -664
rect 1520 -695 1527 -693
rect 1351 -702 1364 -699
rect 927 -709 936 -703
rect 951 -704 1364 -702
rect 927 -726 935 -709
rect 951 -711 994 -704
rect 951 -729 958 -711
rect 1008 -711 1364 -704
rect 1351 -746 1364 -711
rect 1447 -718 1487 -713
rect 1443 -719 1487 -718
rect 490 -842 496 -809
rect 514 -842 521 -798
rect 557 -819 654 -805
rect 557 -820 671 -819
rect 558 -857 755 -839
rect 474 -913 478 -882
rect 558 -898 570 -857
rect 833 -839 845 -837
rect 801 -857 845 -839
rect 915 -838 919 -769
rect 923 -795 1053 -794
rect 932 -804 1053 -795
rect 932 -805 1095 -804
rect 1351 -809 1362 -746
rect 1473 -765 1486 -719
rect 1520 -773 1527 -707
rect 1351 -810 1510 -809
rect 1522 -810 1534 -809
rect 1632 -810 1660 -682
rect 1089 -818 1118 -810
rect 833 -861 845 -857
rect 494 -902 570 -898
rect 558 -903 570 -902
rect 832 -930 845 -861
rect 995 -858 1004 -847
rect 1093 -864 1106 -818
rect 1351 -827 1660 -810
rect 1493 -828 1660 -827
rect 1919 -684 1920 -682
rect 1092 -868 1106 -864
rect 1092 -905 1105 -868
rect 1522 -884 1534 -828
rect 1486 -892 1534 -884
rect 945 -921 1026 -914
rect 832 -932 968 -930
rect 1092 -932 1104 -905
rect 832 -952 1104 -932
rect 985 -1030 1026 -1005
rect 1037 -1030 1039 -1005
rect 1919 -1413 1953 -684
rect 1020 -1414 1958 -1413
rect 1041 -1440 1958 -1414
rect 1919 -1442 1953 -1440
<< m3contact >>
rect 1195 20 1211 32
rect 150 -63 165 -51
rect 588 -110 596 -98
rect 959 -108 985 -95
rect 648 -161 665 -149
rect 479 -223 502 -203
rect 1371 -171 1379 -165
rect 1119 -287 1136 -275
rect 1022 -360 1032 -349
rect 261 -455 295 -430
rect 591 -461 609 -447
rect 1022 -444 1038 -428
rect 591 -598 615 -583
rect 1309 -654 1327 -645
rect 212 -670 227 -659
rect 130 -705 140 -697
rect 260 -787 299 -778
rect 350 -819 366 -811
rect 210 -858 225 -847
rect 488 -809 498 -790
rect 555 -688 565 -683
rect 924 -703 940 -690
rect 994 -713 1008 -704
rect 654 -819 671 -803
rect 755 -862 801 -837
rect 1053 -804 1095 -793
rect 1118 -818 1140 -810
rect 995 -847 1009 -838
rect 1026 -922 1038 -914
rect 413 -1041 426 -1014
rect 1026 -1030 1037 -1002
<< metal3 >>
rect 1196 -26 1210 20
rect 55 -51 63 -50
rect 53 -63 150 -51
rect 55 -124 63 -63
rect 525 -99 535 -98
rect 524 -110 588 -99
rect 958 -108 959 -97
rect 54 -138 63 -124
rect 54 -256 62 -138
rect 525 -176 535 -110
rect 482 -203 498 -202
rect 54 -277 63 -256
rect 55 -322 63 -277
rect 54 -344 63 -322
rect 54 -636 62 -344
rect 260 -455 261 -439
rect 129 -636 136 -635
rect 54 -646 136 -636
rect 129 -697 136 -646
rect 260 -638 295 -455
rect 210 -670 212 -659
rect 129 -702 130 -697
rect 210 -847 223 -670
rect 260 -722 296 -638
rect 482 -690 498 -223
rect 525 -240 536 -176
rect 648 -192 665 -161
rect 648 -204 666 -192
rect 649 -209 666 -204
rect 648 -226 666 -209
rect 525 -451 537 -240
rect 648 -285 665 -226
rect 648 -293 667 -285
rect 650 -361 667 -293
rect 650 -369 668 -361
rect 651 -418 668 -369
rect 650 -445 668 -418
rect 913 -437 932 -144
rect 958 -282 985 -108
rect 1196 -156 1211 -26
rect 1197 -166 1211 -156
rect 1197 -167 1371 -166
rect 1198 -171 1371 -167
rect 960 -403 985 -282
rect 1118 -287 1119 -275
rect 1136 -287 1137 -275
rect 960 -426 986 -403
rect 524 -477 537 -451
rect 591 -447 610 -446
rect 609 -461 610 -447
rect 524 -540 536 -477
rect 523 -584 536 -540
rect 591 -583 610 -461
rect 650 -476 667 -445
rect 650 -502 668 -476
rect 913 -484 933 -437
rect 523 -669 535 -584
rect 523 -673 563 -669
rect 555 -683 562 -673
rect 261 -778 296 -722
rect 261 -790 296 -787
rect 481 -790 501 -690
rect 651 -693 668 -502
rect 914 -690 933 -484
rect 961 -632 986 -426
rect 1022 -428 1031 -360
rect 1118 -406 1137 -287
rect 1117 -476 1137 -406
rect 1117 -490 1139 -476
rect 1119 -543 1139 -490
rect 1118 -560 1139 -543
rect 961 -642 1096 -632
rect 651 -697 669 -693
rect 652 -741 669 -697
rect 914 -702 924 -690
rect 924 -705 933 -703
rect 995 -704 1009 -702
rect 1008 -713 1009 -704
rect 652 -777 670 -741
rect 481 -805 488 -790
rect 498 -805 501 -790
rect 653 -801 670 -777
rect 650 -803 672 -801
rect 650 -819 654 -803
rect 671 -819 672 -803
rect 351 -1056 365 -819
rect 650 -933 672 -819
rect 995 -838 1009 -713
rect 1054 -793 1095 -642
rect 1054 -805 1095 -804
rect 1118 -810 1138 -560
rect 1309 -645 1326 -171
rect 1118 -819 1138 -818
rect 650 -969 674 -933
rect 426 -1015 557 -1014
rect 652 -1015 674 -969
rect 426 -1041 674 -1015
rect 530 -1042 674 -1041
rect 755 -1055 799 -862
rect 1028 -964 1036 -922
rect 1027 -1002 1037 -964
rect 1026 -1031 1037 -1030
rect 394 -1056 803 -1055
rect 351 -1088 803 -1056
rect 351 -1089 760 -1088
use q1c_4_INPUT_OR  q1c_4_INPUT_OR_1
timestamp 1699085113
transform 0 1 1002 -1 0 -1364
box -38 -91 102 31
use q1b_5_INPUT_AND  q1b_5_INPUT_AND_1
timestamp 1699075298
transform 0 1 114 -1 0 -848
box -24 -57 84 37
use 4_input_AND  4_input_AND_2
timestamp 1699820036
transform 0 1 510 -1 0 -920
box -22 -53 85 30
use q1a_NOT  q1a_NOT_7
timestamp 1698924755
transform 0 1 491 -1 0 -859
box -12 -23 15 29
use 3_input_AND  3_input_AND_1
timestamp 1699847323
transform 0 1 944 -1 0 -840
box -19 -42 67 25
use 2_input_AND  2_input_AND_1
timestamp 1699478438
transform 0 1 1449 -1 0 -931
box -12 -30 69 33
use q1a_NOT  q1a_NOT_6
timestamp 1698924755
transform 0 1 79 -1 0 -730
box -12 -23 15 29
use q1a_NOT  q1a_NOT_5
timestamp 1698924755
transform 0 1 928 -1 0 -743
box -12 -23 15 29
use q1c_4_INPUT_OR  q1c_4_INPUT_OR_0
timestamp 1699085113
transform 1 0 1602 0 1 -387
box -38 -91 102 31
use q1a_NOT  q1a_NOT_4
timestamp 1698924755
transform 0 1 1442 -1 0 -685
box -12 -23 15 29
use q1b_5_INPUT_AND  q1b_5_INPUT_AND_0
timestamp 1699075298
transform 0 1 174 -1 0 -185
box -24 -57 84 37
use q1a_NOT  q1a_NOT_3
timestamp 1698924755
transform 0 1 158 -1 0 -123
box -12 -23 15 29
use 4_input_AND  4_input_AND_1
timestamp 1699820036
transform 0 1 606 -1 0 -205
box -22 -53 85 30
use q1a_NOT  q1a_NOT_2
timestamp 1698924755
transform 0 1 591 -1 0 -130
box -12 -23 15 29
use 3_input_AND  3_input_AND_0
timestamp 1699847323
transform 0 1 1031 -1 0 -194
box -19 -42 67 25
use q1a_NOT  q1a_NOT_1
timestamp 1698924755
transform 0 1 1015 -1 0 -129
box -12 -23 15 29
use 2_input_AND  2_input_AND_0
timestamp 1699478438
transform 0 1 1418 -1 0 -186
box -12 -30 69 33
use q1a_NOT  q1a_NOT_0
timestamp 1698924755
transform 0 1 1413 -1 0 -138
box -12 -23 15 29
use XNOR  XNOR_0
timestamp 1699711768
transform 1 0 19 0 1 17
box -19 -17 270 145
use XNOR  XNOR_1
timestamp 1699711768
transform 1 0 447 0 1 17
box -19 -17 270 145
use XNOR  XNOR_2
timestamp 1699711768
transform 1 0 869 0 1 16
box -19 -17 270 145
use XNOR  XNOR_3
timestamp 1699711768
transform 1 0 1268 0 1 23
box -19 -17 270 145
use 4_input_AND  4_input_AND_0
timestamp 1699820036
transform 1 0 1624 0 1 100
box -22 -53 85 30
<< labels >>
rlabel metal1 -2 1 1 4 1 GND
rlabel metal1 -4 88 -2 90 1 A0
rlabel metal1 161 8 163 9 1 B0
rlabel metal1 286 93 287 94 1 A0B0
rlabel metal1 425 89 426 90 1 A1
rlabel metal1 587 8 588 9 1 B1
rlabel metal1 714 93 715 94 1 A1B1
rlabel metal1 847 88 848 89 1 A2
rlabel metal1 1011 7 1012 8 1 B2
rlabel metal1 1139 92 1140 93 1 A2B2
rlabel metal1 1245 95 1246 96 1 A3
rlabel metal1 1411 14 1412 15 1 B3
rlabel metal1 1535 99 1537 100 1 A3B3
rlabel metal1 -22 144 -20 145 3 VDD
rlabel metal1 1708 95 1709 96 1 A_IS_EQUAL_B
rlabel metal1 592 -147 593 -146 1 B1_NOT
rlabel metal1 1015 -149 1016 -147 1 B2_NOT
rlabel metal1 1414 -156 1415 -155 1 B3_NOT
rlabel metal1 159 -139 160 -138 1 B0_NOT
rlabel metal1 1420 -258 1421 -257 1 A3_B3NOT
rlabel metal1 1026 -265 1027 -264 1 A2_B2NOT_A3B3XNOR
rlabel metal1 1712 -408 1714 -406 1 A_greater_than_B
rlabel metal1 179 -271 180 -270 1 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR
rlabel metal1 602 -287 604 -286 1 A1_B1NOT_A3B3XNOR_A2B2XOR
rlabel metal1 928 -759 930 -757 1 A2NOT
rlabel m2contact 80 -746 81 -743 1 A0NOT
rlabel metal1 492 -878 494 -876 1 A1NOT
rlabel metal1 1450 -1002 1452 -1001 1 A3NOT_B3
rlabel metal1 939 -910 940 -908 1 A2NOT_B2_A3B3XNOR
rlabel metal1 505 -1002 506 -1000 1 A1NOTB1_A2XNORB2_A3XNORB3
rlabel metal1 119 -935 121 -934 1 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3
rlabel metal1 980 -1472 983 -1468 1 A_less_than_B
<< end >>
