.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include decoder.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'
V_in_S0 node_S0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_S1 node_S1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)

* V_in_S1 node_S1 gnd DC 1.8
* V_in_S0 node_S0 gnd DC 0

X1 node_S0 node_S1 node_D0 node_D1 node_D2 node_D3 node_x gnd decoder

C1 node_out gnd 100f

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_S0) v(node_S1)+2 v(node_D0)+4 v(node_D1)+6 v(node_D2)+8 v(node_D3)+10
* plot v(node_D0) v(node_D1)+2 v(node_D2)+4 v(node_D3)+6
.end
.endc
