magic
tech scmos
timestamp 1699820036
<< nwell >>
rect -22 4 30 23
rect 40 5 75 21
<< ntransistor >>
rect 56 -28 58 -24
rect -10 -45 -8 -38
rect -1 -45 1 -38
rect 8 -45 10 -38
rect 17 -45 19 -38
<< ptransistor >>
rect -10 11 -8 17
rect -1 11 1 17
rect 8 11 10 17
rect 17 11 19 17
rect 56 11 58 15
<< ndiffusion >>
rect 53 -28 56 -24
rect 58 -28 62 -24
rect -11 -45 -10 -38
rect -8 -45 -1 -38
rect 1 -45 8 -38
rect 10 -45 17 -38
rect 19 -45 22 -38
<< pdiffusion >>
rect -11 11 -10 17
rect -8 11 -7 17
rect -3 11 -1 17
rect 1 11 2 17
rect 6 11 8 17
rect 10 11 12 17
rect 16 11 17 17
rect 19 11 20 17
rect 53 11 56 15
rect 58 11 62 15
<< ndcontact >>
rect 49 -28 53 -24
rect 62 -28 66 -24
rect -15 -45 -11 -38
rect 22 -45 26 -38
<< pdcontact >>
rect -15 11 -11 17
rect -7 11 -3 17
rect 2 11 6 17
rect 12 11 16 17
rect 20 11 24 17
rect 49 11 53 15
rect 62 11 66 15
<< polysilicon >>
rect -10 17 -8 20
rect -1 17 1 20
rect 8 17 10 21
rect 17 17 19 20
rect 56 15 58 19
rect -10 -12 -8 11
rect -10 -38 -8 -16
rect -1 -18 1 11
rect -1 -38 1 -22
rect 8 -25 10 11
rect 8 -38 10 -29
rect 17 -32 19 11
rect 56 -2 58 11
rect 57 -7 58 -2
rect 56 -24 58 -7
rect 17 -38 19 -36
rect -10 -50 -8 -45
rect -1 -49 1 -45
rect 8 -49 10 -45
rect 17 -49 19 -45
rect 56 -50 58 -28
<< polycontact >>
rect -12 -16 -8 -12
rect -3 -22 1 -18
rect 6 -29 10 -25
rect 52 -7 57 -2
rect 15 -36 19 -32
<< metal1 >>
rect -22 25 83 30
rect -7 17 -3 25
rect 12 17 16 25
rect 49 15 53 25
rect -15 -2 -11 11
rect 2 -2 6 11
rect 20 -2 24 11
rect 62 -2 66 11
rect -15 -7 52 -2
rect 62 -7 76 -2
rect -14 -16 -12 -12
rect -5 -22 -3 -18
rect 4 -29 6 -25
rect 13 -36 15 -32
rect 22 -38 26 -7
rect 62 -24 66 -7
rect -15 -48 -11 -45
rect 49 -48 53 -28
rect -19 -53 85 -48
<< labels >>
rlabel metal1 29 27 31 28 5 VDD
rlabel metal1 71 -6 72 -5 1 OUT_FINAL
rlabel metal1 44 -5 45 -4 1 OUT
rlabel metal1 14 -34 15 -33 1 D
rlabel metal1 5 -27 6 -26 1 C
rlabel metal1 -4 -21 -3 -20 1 B
rlabel metal1 -13 -14 -12 -13 1 A
rlabel metal1 38 -51 39 -50 1 GND
<< end >>
