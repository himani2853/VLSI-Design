magic
tech scmos
timestamp 1699075298
<< nwell >>
rect -24 8 40 29
rect 50 10 82 29
<< ntransistor >>
rect 65 -10 67 -4
rect -13 -43 -11 -36
rect -3 -43 -1 -36
rect 6 -43 8 -36
rect 15 -43 17 -36
rect 24 -43 26 -36
<< ptransistor >>
rect -13 14 -11 21
rect -3 14 -1 21
rect 6 14 8 21
rect 15 14 17 21
rect 24 14 26 21
rect 65 17 67 23
<< ndiffusion >>
rect 63 -10 65 -4
rect 67 -10 70 -4
rect -15 -43 -13 -36
rect -11 -43 -3 -36
rect -1 -43 6 -36
rect 8 -43 15 -36
rect 17 -43 24 -36
rect 26 -43 29 -36
<< pdiffusion >>
rect -14 14 -13 21
rect -11 14 -8 21
rect -4 14 -3 21
rect -1 14 1 21
rect 5 14 6 21
rect 8 14 9 21
rect 13 14 15 21
rect 17 14 18 21
rect 22 14 24 21
rect 26 14 29 21
rect 63 17 65 23
rect 67 17 70 23
<< ndcontact >>
rect 57 -10 63 -4
rect 70 -10 75 -4
rect -19 -43 -15 -36
rect 29 -43 33 -36
<< pdcontact >>
rect -18 14 -14 21
rect -8 14 -4 21
rect 1 14 5 21
rect 9 14 13 21
rect 18 14 22 21
rect 29 14 33 21
rect 57 17 63 23
rect 70 17 75 23
<< polysilicon >>
rect -13 21 -11 25
rect -3 21 -1 25
rect 6 21 8 25
rect 15 21 17 25
rect 24 21 26 25
rect 65 23 67 26
rect -13 8 -11 14
rect -13 -36 -11 4
rect -3 0 -1 14
rect -3 -36 -1 -4
rect 6 -8 8 14
rect 6 -36 8 -12
rect 15 -16 17 14
rect 15 -36 17 -20
rect 24 -24 26 14
rect 65 7 67 17
rect 65 -4 67 3
rect 65 -14 67 -10
rect 24 -36 26 -28
rect -13 -47 -11 -43
rect -3 -47 -1 -43
rect 6 -47 8 -43
rect 15 -47 17 -43
rect 24 -47 26 -43
<< polycontact >>
rect -16 4 -11 8
rect -7 -4 -1 0
rect 3 -12 8 -8
rect 13 -20 18 -16
rect 53 3 67 7
rect 21 -28 26 -24
<< metal1 >>
rect -24 29 82 37
rect -18 21 -14 29
rect 1 21 5 29
rect 18 21 22 29
rect 57 23 63 29
rect -20 4 -16 8
rect -8 7 -4 14
rect 9 7 13 14
rect 29 7 33 14
rect 70 7 75 17
rect -8 3 53 7
rect 70 3 84 7
rect -20 -4 -7 0
rect -20 -12 3 -8
rect -20 -20 13 -16
rect -20 -28 21 -24
rect 29 -36 33 3
rect 70 -4 75 3
rect 57 -15 63 -10
rect 57 -20 83 -15
rect -19 -49 -15 -43
rect 78 -49 83 -20
rect -19 -57 83 -49
<< labels >>
rlabel metal1 2 34 12 36 5 VDD
rlabel metal1 43 3 53 5 1 OUT
rlabel metal1 -18 4 -16 6 1 A
rlabel metal1 -17 -4 -15 -2 1 B
rlabel metal1 -17 -12 -15 -10 1 C
rlabel metal1 -17 -20 -15 -18 1 D
rlabel metal1 -17 -28 -15 -26 1 E
rlabel metal1 3 -57 9 -53 1 GND
rlabel metal1 79 5 83 7 7 OUT_FINAL
<< end >>
