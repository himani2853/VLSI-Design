* SPICE3 file created from q1a_NOT.ext - technology: scmos
.include TSMC_180nm.txt


.param SUPPLY = 1.8


.global GND

Vdd VDD GND 'SUPPLY'

V_in_in in GND PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
.option scale=0.09u

M1000 out in vdd VDD CMOSP w=6 l=2
+  ad=36 pd=24 as=30 ps=22
M1001 out in gnd Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=30 ps=22
C0 vdd VDD 0.05fF
C1 in gnd 0.04fF
C2 in VDD 0.07fF
C3 out vdd 0.10fF
C4 out gnd 0.10fF
C5 out in 0.04fF
C6 out VDD 0.04fF
C7 gnd Gnd 0.11fF
C8 out Gnd 0.06fF
C9 vdd Gnd 0.06fF
C10 in Gnd 0.14fF
C11 VDD Gnd 0.50fF
.tran 1n 500n

.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(in) v(out)+2
* plot v(OUT_FINAL)/
* hardcopy image.ps v(node_a) v(node_b)+2 v(OUT)+4
.end
.endc