* SPICE3 file created from alu_complete.ext - technology: scmos
.include TSMC_180nm.txt



.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}

.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}


.param wp1 = wn1
.param wp2 = wn1

.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}


.global GND

* 1010-10
* 1001-9
* 0110
* 0111
* 0001
* 10011
Vdd VDD GND 'SUPPLY'
V_in_S0_DECODER S0_DECODER GND DC 1.8
V_in_S1_DECODER S1_DECODER GND DC 1.8

V_in_INPUT_ALU_A0 INPUT_ALU_A0 GND PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_INPUT_ALU_A1 INPUT_ALU_A1 GND PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_INPUT_ALU_A2 INPUT_ALU_A2 GND PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_INPUT_ALU_A3 INPUT_ALU_A3 GND PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
* 0110
* 1101
* 10011
* V_in_M M gnd DC 1.8
V_in_INPUT_ALU_B0 INPUT_ALU_B0 GND DC 1.8
V_in_INPUT_ALU_B1 INPUT_ALU_B1 GND DC 1.8
V_in_INPUT_ALU_B2 INPUT_ALU_B2 GND DC 1.8
V_in_INPUT_ALU_B3 INPUT_ALU_B3 GND DC 1.8
.option scale=0.09u


M1000 VDD OUTPUT_ALU_ANDBLOCK_B0 and_block_0/2_input_AND_0/OUT and_block_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=6526 pd=4768 as=24 ps=20
M1001 and_block_0/2_input_AND_0/a_4_n21# OUTPUT_ALU_ANDBLOCK_A0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=5033 ps=3668
M1002 AND_OUTPUT_A0B0 and_block_0/2_input_AND_0/OUT VDD and_block_0/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1003 and_block_0/2_input_AND_0/OUT OUTPUT_ALU_ANDBLOCK_A0 VDD and_block_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 AND_OUTPUT_A0B0 and_block_0/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 and_block_0/2_input_AND_0/OUT OUTPUT_ALU_ANDBLOCK_B0 and_block_0/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1006 VDD OUTPUT_ALU_ANDBLOCK_B1 and_block_0/2_input_AND_1/OUT and_block_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1007 and_block_0/2_input_AND_1/a_4_n21# OUTPUT_ALU_ANDBLOCK_A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1008 AND_OUTPUT_A1B1 and_block_0/2_input_AND_1/OUT VDD and_block_0/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1009 and_block_0/2_input_AND_1/OUT OUTPUT_ALU_ANDBLOCK_A1 VDD and_block_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 AND_OUTPUT_A1B1 and_block_0/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1011 and_block_0/2_input_AND_1/OUT OUTPUT_ALU_ANDBLOCK_B1 and_block_0/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1012 VDD OUTPUT_ALU_ANDBLOCK_B2 and_block_0/2_input_AND_2/OUT and_block_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1013 and_block_0/2_input_AND_2/a_4_n21# OUTPUT_ALU_ANDBLOCK_A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1014 AND_OUTPUT_A2B2 and_block_0/2_input_AND_2/OUT VDD and_block_0/2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1015 and_block_0/2_input_AND_2/OUT OUTPUT_ALU_ANDBLOCK_A2 VDD and_block_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 AND_OUTPUT_A2B2 and_block_0/2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1017 and_block_0/2_input_AND_2/OUT OUTPUT_ALU_ANDBLOCK_B2 and_block_0/2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1018 VDD OUTPUT_ALU_ANDBLOCK_B3 and_block_0/2_input_AND_3/OUT and_block_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1019 and_block_0/2_input_AND_3/a_4_n21# OUTPUT_ALU_ANDBLOCK_A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1020 AND_OUTPUT_A3B3 and_block_0/2_input_AND_3/OUT VDD and_block_0/2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1021 and_block_0/2_input_AND_3/OUT OUTPUT_ALU_ANDBLOCK_A3 VDD and_block_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 AND_OUTPUT_A3B3 and_block_0/2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1023 and_block_0/2_input_AND_3/OUT OUTPUT_ALU_ANDBLOCK_B3 and_block_0/2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1024 VDD adder_subtractor_0/B0_XOR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1025 adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=76 pd=62 as=44 ps=38
M1026 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/B0_XOR GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 VDD OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/B0_XOR OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=48 ps=40
M1029 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_A0 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1030 adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A0 Gnd CMOSN w=4 l=3
+  ad=72 pd=60 as=48 ps=40
M1031 adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/B0_XOR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1032 VDD ADD_SUB_M adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1033 ADDER_SUB_S0 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1034 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1035 VDD adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 ADDER_SUB_S0 ADD_SUB_M adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1037 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_0/AXORB GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1038 ADDER_SUB_S0 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_0/AXORB Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1039 ADDER_SUB_S0 ADD_SUB_M adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1040 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT adder_subtractor_0/full_adder_0/2_input_OR_0/A GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1041 adder_subtractor_0/full_adder_0/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_0/2_input_OR_0/A VDD adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1042 ADDER_SUB_C1 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT VDD adder_subtractor_0/full_adder_0/2_input_OR_0/w_30_15# CMOSP w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1043 ADDER_SUB_C1 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1044 GND adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1046 VDD OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1047 adder_subtractor_0/full_adder_0/2_input_AND_0/a_4_n21# adder_subtractor_0/B0_XOR GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1048 adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_AND_0/OUT VDD adder_subtractor_0/full_adder_0/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1049 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT adder_subtractor_0/B0_XOR VDD adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1051 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1052 VDD adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/2_input_AND_1/OUT adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1053 adder_subtractor_0/full_adder_0/2_input_AND_1/a_4_n21# ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1054 adder_subtractor_0/full_adder_0/2_input_OR_0/A adder_subtractor_0/full_adder_0/2_input_AND_1/OUT VDD adder_subtractor_0/full_adder_0/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1055 adder_subtractor_0/full_adder_0/2_input_AND_1/OUT ADD_SUB_M VDD adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 adder_subtractor_0/full_adder_0/2_input_OR_0/A adder_subtractor_0/full_adder_0/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1057 adder_subtractor_0/full_adder_0/2_input_AND_1/OUT adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1058 VDD OUTPUT_ALU_ADDER_A1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1059 adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=76 pd=62 as=44 ps=38
M1060 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1061 VDD adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 adder_subtractor_0/full_adder_1/AXORB OUTPUT_ALU_ADDER_A1 adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=76 ps=62
M1063 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B1_XOR GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1064 adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/B1_XOR Gnd CMOSN w=4 l=3
+  ad=72 pd=60 as=72 ps=60
M1065 adder_subtractor_0/full_adder_1/AXORB OUTPUT_ALU_ADDER_A1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1066 VDD ADDER_SUB_C1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1067 ADDER_SUB_S1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1068 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1069 VDD adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1070 ADDER_SUB_S1 ADDER_SUB_C1 adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1071 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_1/AXORB GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1072 ADDER_SUB_S1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_1/AXORB Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1073 ADDER_SUB_S1 ADDER_SUB_C1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1074 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT adder_subtractor_0/full_adder_1/2_input_OR_0/A GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1075 adder_subtractor_0/full_adder_1/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_1/2_input_OR_0/A VDD adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1076 ADDER_SUB_C2 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT VDD adder_subtractor_0/full_adder_1/2_input_OR_0/w_30_15# CMOSP w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1077 ADDER_SUB_C2 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1078 GND adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1080 VDD adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/2_input_AND_0/OUT adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1081 adder_subtractor_0/full_adder_1/2_input_AND_0/a_4_n21# OUTPUT_ALU_ADDER_A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1082 adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_AND_0/OUT VDD adder_subtractor_0/full_adder_1/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1083 adder_subtractor_0/full_adder_1/2_input_AND_0/OUT OUTPUT_ALU_ADDER_A1 VDD adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1085 adder_subtractor_0/full_adder_1/2_input_AND_0/OUT adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1086 VDD adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/2_input_AND_1/OUT adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1087 adder_subtractor_0/full_adder_1/2_input_AND_1/a_4_n21# ADDER_SUB_C1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1088 adder_subtractor_0/full_adder_1/2_input_OR_0/A adder_subtractor_0/full_adder_1/2_input_AND_1/OUT VDD adder_subtractor_0/full_adder_1/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1089 adder_subtractor_0/full_adder_1/2_input_AND_1/OUT ADDER_SUB_C1 VDD adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 adder_subtractor_0/full_adder_1/2_input_OR_0/A adder_subtractor_0/full_adder_1/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1091 adder_subtractor_0/full_adder_1/2_input_AND_1/OUT adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1092 VDD OUTPUT_ALU_ADDER_B0 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1093 adder_subtractor_0/B0_XOR adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1094 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_B0 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1095 VDD ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 adder_subtractor_0/B0_XOR OUTPUT_ALU_ADDER_B0 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=120 ps=100
M1097 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1098 adder_subtractor_0/B0_XOR adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR ADD_SUB_M Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=120 ps=100
M1099 adder_subtractor_0/B0_XOR OUTPUT_ALU_ADDER_B0 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1100 VDD OUTPUT_ALU_ADDER_A2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1101 adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=76 pd=62 as=44 ps=38
M1102 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1103 VDD adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 adder_subtractor_0/full_adder_2/AXORB OUTPUT_ALU_ADDER_A2 adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=76 ps=62
M1105 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B2_XOR GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1106 adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/B2_XOR Gnd CMOSN w=4 l=3
+  ad=72 pd=60 as=72 ps=60
M1107 adder_subtractor_0/full_adder_2/AXORB OUTPUT_ALU_ADDER_A2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1108 VDD ADDER_SUB_C2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1109 ADDER_SUB_S2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1110 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1111 VDD adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 ADDER_SUB_S2 ADDER_SUB_C2 adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1113 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_2/AXORB GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1114 ADDER_SUB_S2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_2/AXORB Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1115 ADDER_SUB_S2 ADDER_SUB_C2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1116 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT adder_subtractor_0/full_adder_2/2_input_OR_0/A GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1117 adder_subtractor_0/full_adder_2/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_2/2_input_OR_0/A VDD adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1118 ADDER_SUB_C3 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT VDD adder_subtractor_0/full_adder_2/2_input_OR_0/w_30_15# CMOSP w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1119 ADDER_SUB_C3 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1120 GND adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1122 VDD adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/2_input_AND_0/OUT adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1123 adder_subtractor_0/full_adder_2/2_input_AND_0/a_4_n21# OUTPUT_ALU_ADDER_A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1124 adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_AND_0/OUT VDD adder_subtractor_0/full_adder_2/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1125 adder_subtractor_0/full_adder_2/2_input_AND_0/OUT OUTPUT_ALU_ADDER_A2 VDD adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1127 adder_subtractor_0/full_adder_2/2_input_AND_0/OUT adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1128 VDD adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/2_input_AND_1/OUT adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1129 adder_subtractor_0/full_adder_2/2_input_AND_1/a_4_n21# ADDER_SUB_C2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1130 adder_subtractor_0/full_adder_2/2_input_OR_0/A adder_subtractor_0/full_adder_2/2_input_AND_1/OUT VDD adder_subtractor_0/full_adder_2/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1131 adder_subtractor_0/full_adder_2/2_input_AND_1/OUT ADDER_SUB_C2 VDD adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 adder_subtractor_0/full_adder_2/2_input_OR_0/A adder_subtractor_0/full_adder_2/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1133 adder_subtractor_0/full_adder_2/2_input_AND_1/OUT adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1134 VDD OUTPUT_ALU_ADDER_A3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1135 adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=76 pd=62 as=44 ps=38
M1136 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1137 VDD adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1138 adder_subtractor_0/full_adder_3/AXORB OUTPUT_ALU_ADDER_A3 adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=76 ps=62
M1139 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B3_XOR GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1140 adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/B3_XOR Gnd CMOSN w=4 l=3
+  ad=72 pd=60 as=72 ps=60
M1141 adder_subtractor_0/full_adder_3/AXORB OUTPUT_ALU_ADDER_A3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1142 VDD ADDER_SUB_C3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1143 ADDER_SUB_S3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1144 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1145 VDD adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 ADDER_SUB_S3 ADDER_SUB_C3 adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1147 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_3/AXORB GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1148 ADDER_SUB_S3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/full_adder_3/AXORB Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1149 ADDER_SUB_S3 ADDER_SUB_C3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1150 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT adder_subtractor_0/full_adder_3/2_input_OR_0/A GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1151 adder_subtractor_0/full_adder_3/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_3/2_input_OR_0/A VDD adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1152 ADDER_SUB_C4 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT VDD adder_subtractor_0/full_adder_3/2_input_OR_0/w_30_15# CMOSP w=5 l=2
+  ad=64 pd=46 as=0 ps=0
M1153 ADDER_SUB_C4 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=64 pd=46 as=0 ps=0
M1154 GND adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_OR_0/a_n7_22# adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1156 VDD adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/2_input_AND_0/OUT adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1157 adder_subtractor_0/full_adder_3/2_input_AND_0/a_4_n21# OUTPUT_ALU_ADDER_A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1158 adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_AND_0/OUT VDD adder_subtractor_0/full_adder_3/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1159 adder_subtractor_0/full_adder_3/2_input_AND_0/OUT OUTPUT_ALU_ADDER_A3 VDD adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1161 adder_subtractor_0/full_adder_3/2_input_AND_0/OUT adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1162 VDD adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/2_input_AND_1/OUT adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1163 adder_subtractor_0/full_adder_3/2_input_AND_1/a_4_n21# ADDER_SUB_C3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1164 adder_subtractor_0/full_adder_3/2_input_OR_0/A adder_subtractor_0/full_adder_3/2_input_AND_1/OUT VDD adder_subtractor_0/full_adder_3/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1165 adder_subtractor_0/full_adder_3/2_input_AND_1/OUT ADDER_SUB_C3 VDD adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 adder_subtractor_0/full_adder_3/2_input_OR_0/A adder_subtractor_0/full_adder_3/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1167 adder_subtractor_0/full_adder_3/2_input_AND_1/OUT adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1168 VDD OUTPUT_ALU_ADDER_B1 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1169 adder_subtractor_0/B1_XOR adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_53_n17# CMOSP w=4 l=3
+  ad=0 pd=0 as=44 ps=38
M1170 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR OUTPUT_ALU_ADDER_B1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1171 VDD ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1172 adder_subtractor_0/B1_XOR OUTPUT_ALU_ADDER_B1 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1173 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1174 adder_subtractor_0/B1_XOR adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR ADD_SUB_M Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1175 adder_subtractor_0/B1_XOR OUTPUT_ALU_ADDER_B1 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1176 VDD OUTPUT_ALU_ADDER_B2 adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_2/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1177 adder_subtractor_0/B2_XOR adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_2/w_53_n17# CMOSP w=4 l=3
+  ad=0 pd=0 as=44 ps=38
M1178 adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR OUTPUT_ALU_ADDER_B2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1179 VDD ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_2/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 adder_subtractor_0/B2_XOR OUTPUT_ALU_ADDER_B2 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1181 adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1182 adder_subtractor_0/B2_XOR adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR ADD_SUB_M Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1183 adder_subtractor_0/B2_XOR OUTPUT_ALU_ADDER_B2 adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1184 VDD OUTPUT_ALU_ADDER_B3 adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_3/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1185 adder_subtractor_0/B3_XOR adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_3/w_53_n17# CMOSP w=4 l=3
+  ad=0 pd=0 as=44 ps=38
M1186 adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR OUTPUT_ALU_ADDER_B3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1187 VDD ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_3/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 adder_subtractor_0/B3_XOR OUTPUT_ALU_ADDER_B3 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1189 adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1190 adder_subtractor_0/B3_XOR adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR ADD_SUB_M Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1191 adder_subtractor_0/B3_XOR OUTPUT_ALU_ADDER_B3 adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1192 VDD ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_4/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1193 ADDER_SUB_CFINAL adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_4/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1194 adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1195 VDD ADDER_SUB_C4 adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_4/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 ADDER_SUB_CFINAL ADD_SUB_M ADDER_SUB_C4 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1197 adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR ADDER_SUB_C4 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1198 ADDER_SUB_CFINAL adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR ADDER_SUB_C4 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1199 ADDER_SUB_CFINAL ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1200 VDD S0_S1_DECODER enable_0/2_input_AND_7/OUT enable_0/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1201 enable_0/2_input_AND_7/a_4_n21# INPUT_ALU_B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1202 OUTPUT_ALU_ANDBLOCK_B3 enable_0/2_input_AND_7/OUT VDD enable_0/2_input_AND_7/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1203 enable_0/2_input_AND_7/OUT INPUT_ALU_B3 VDD enable_0/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 OUTPUT_ALU_ANDBLOCK_B3 enable_0/2_input_AND_7/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1205 enable_0/2_input_AND_7/OUT S0_S1_DECODER enable_0/2_input_AND_7/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1206 VDD S0_S1_DECODER enable_0/2_input_AND_0/OUT enable_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1207 enable_0/2_input_AND_0/a_4_n21# INPUT_ALU_A0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1208 OUTPUT_ALU_ANDBLOCK_A0 enable_0/2_input_AND_0/OUT VDD enable_0/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1209 enable_0/2_input_AND_0/OUT INPUT_ALU_A0 VDD enable_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1210 OUTPUT_ALU_ANDBLOCK_A0 enable_0/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1211 enable_0/2_input_AND_0/OUT S0_S1_DECODER enable_0/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1212 VDD S0_S1_DECODER enable_0/2_input_AND_1/OUT enable_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1213 enable_0/2_input_AND_1/a_4_n21# INPUT_ALU_A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1214 OUTPUT_ALU_ANDBLOCK_A1 enable_0/2_input_AND_1/OUT VDD enable_0/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1215 enable_0/2_input_AND_1/OUT INPUT_ALU_A1 VDD enable_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 OUTPUT_ALU_ANDBLOCK_A1 enable_0/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1217 enable_0/2_input_AND_1/OUT S0_S1_DECODER enable_0/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1218 VDD S0_S1_DECODER enable_0/2_input_AND_2/OUT enable_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1219 enable_0/2_input_AND_2/a_4_n21# INPUT_ALU_A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1220 OUTPUT_ALU_ANDBLOCK_A2 enable_0/2_input_AND_2/OUT VDD enable_0/2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1221 enable_0/2_input_AND_2/OUT INPUT_ALU_A2 VDD enable_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1222 OUTPUT_ALU_ANDBLOCK_A2 enable_0/2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1223 enable_0/2_input_AND_2/OUT S0_S1_DECODER enable_0/2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1224 VDD S0_S1_DECODER enable_0/2_input_AND_3/OUT enable_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1225 enable_0/2_input_AND_3/a_4_n21# INPUT_ALU_A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1226 OUTPUT_ALU_ANDBLOCK_A3 enable_0/2_input_AND_3/OUT VDD enable_0/2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1227 enable_0/2_input_AND_3/OUT INPUT_ALU_A3 VDD enable_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 OUTPUT_ALU_ANDBLOCK_A3 enable_0/2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1229 enable_0/2_input_AND_3/OUT S0_S1_DECODER enable_0/2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1230 VDD S0_S1_DECODER enable_0/2_input_AND_4/OUT enable_0/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1231 enable_0/2_input_AND_4/a_4_n21# INPUT_ALU_B0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1232 OUTPUT_ALU_ANDBLOCK_B0 enable_0/2_input_AND_4/OUT VDD enable_0/2_input_AND_4/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1233 enable_0/2_input_AND_4/OUT INPUT_ALU_B0 VDD enable_0/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 OUTPUT_ALU_ANDBLOCK_B0 enable_0/2_input_AND_4/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1235 enable_0/2_input_AND_4/OUT S0_S1_DECODER enable_0/2_input_AND_4/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1236 VDD S0_S1_DECODER enable_0/2_input_AND_5/OUT enable_0/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1237 enable_0/2_input_AND_5/a_4_n21# INPUT_ALU_B1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1238 OUTPUT_ALU_ANDBLOCK_B1 enable_0/2_input_AND_5/OUT VDD enable_0/2_input_AND_5/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1239 enable_0/2_input_AND_5/OUT INPUT_ALU_B1 VDD enable_0/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 OUTPUT_ALU_ANDBLOCK_B1 enable_0/2_input_AND_5/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1241 enable_0/2_input_AND_5/OUT S0_S1_DECODER enable_0/2_input_AND_5/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1242 VDD S0_S1_DECODER enable_0/2_input_AND_6/OUT enable_0/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1243 enable_0/2_input_AND_6/a_4_n21# INPUT_ALU_B2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1244 OUTPUT_ALU_ANDBLOCK_B2 enable_0/2_input_AND_6/OUT VDD enable_0/2_input_AND_6/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1245 enable_0/2_input_AND_6/OUT INPUT_ALU_B2 VDD enable_0/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 OUTPUT_ALU_ANDBLOCK_B2 enable_0/2_input_AND_6/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1247 enable_0/2_input_AND_6/OUT S0_S1_DECODER enable_0/2_input_AND_6/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1248 VDD S0BAR_S1_DECODER enable_1/2_input_AND_7/OUT enable_1/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1249 enable_1/2_input_AND_7/a_4_n21# INPUT_ALU_B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1250 OUTPUT_ALU_COMPARATOR_B3 enable_1/2_input_AND_7/OUT VDD enable_1/2_input_AND_7/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1251 enable_1/2_input_AND_7/OUT INPUT_ALU_B3 VDD enable_1/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 OUTPUT_ALU_COMPARATOR_B3 enable_1/2_input_AND_7/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1253 enable_1/2_input_AND_7/OUT S0BAR_S1_DECODER enable_1/2_input_AND_7/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1254 VDD S0BAR_S1_DECODER enable_1/2_input_AND_0/OUT enable_1/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1255 enable_1/2_input_AND_0/a_4_n21# INPUT_ALU_A0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1256 OUTPUT_ALU_COMPARATOR_A0 enable_1/2_input_AND_0/OUT VDD enable_1/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1257 enable_1/2_input_AND_0/OUT INPUT_ALU_A0 VDD enable_1/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 OUTPUT_ALU_COMPARATOR_A0 enable_1/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1259 enable_1/2_input_AND_0/OUT S0BAR_S1_DECODER enable_1/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1260 VDD S0BAR_S1_DECODER enable_1/2_input_AND_1/OUT enable_1/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1261 enable_1/2_input_AND_1/a_4_n21# INPUT_ALU_A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1262 OUTPUT_ALU_COMPARATOR_A1 enable_1/2_input_AND_1/OUT VDD enable_1/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1263 enable_1/2_input_AND_1/OUT INPUT_ALU_A1 VDD enable_1/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 OUTPUT_ALU_COMPARATOR_A1 enable_1/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1265 enable_1/2_input_AND_1/OUT S0BAR_S1_DECODER enable_1/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1266 VDD S0BAR_S1_DECODER enable_1/2_input_AND_2/OUT enable_1/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1267 enable_1/2_input_AND_2/a_4_n21# INPUT_ALU_A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1268 OUTPUT_ALU_COMPARATOR_A2 enable_1/2_input_AND_2/OUT VDD enable_1/2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1269 enable_1/2_input_AND_2/OUT INPUT_ALU_A2 VDD enable_1/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 OUTPUT_ALU_COMPARATOR_A2 enable_1/2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1271 enable_1/2_input_AND_2/OUT S0BAR_S1_DECODER enable_1/2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1272 VDD S0BAR_S1_DECODER enable_1/2_input_AND_3/OUT enable_1/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1273 enable_1/2_input_AND_3/a_4_n21# INPUT_ALU_A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1274 OUTPUT_ALU_COMPARATOR_A3 enable_1/2_input_AND_3/OUT VDD enable_1/2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1275 enable_1/2_input_AND_3/OUT INPUT_ALU_A3 VDD enable_1/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 OUTPUT_ALU_COMPARATOR_A3 enable_1/2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=48 pd=40 as=0 ps=0
M1277 enable_1/2_input_AND_3/OUT S0BAR_S1_DECODER enable_1/2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1278 VDD S0BAR_S1_DECODER enable_1/2_input_AND_4/OUT enable_1/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1279 enable_1/2_input_AND_4/a_4_n21# INPUT_ALU_B0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1280 OUTPUT_ALU_COMPARATOR_B0 enable_1/2_input_AND_4/OUT VDD enable_1/2_input_AND_4/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1281 enable_1/2_input_AND_4/OUT INPUT_ALU_B0 VDD enable_1/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 OUTPUT_ALU_COMPARATOR_B0 enable_1/2_input_AND_4/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1283 enable_1/2_input_AND_4/OUT S0BAR_S1_DECODER enable_1/2_input_AND_4/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1284 VDD S0BAR_S1_DECODER enable_1/2_input_AND_5/OUT enable_1/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1285 enable_1/2_input_AND_5/a_4_n21# INPUT_ALU_B1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1286 OUTPUT_ALU_COMPARATOR_B1 enable_1/2_input_AND_5/OUT VDD enable_1/2_input_AND_5/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1287 enable_1/2_input_AND_5/OUT INPUT_ALU_B1 VDD enable_1/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1288 OUTPUT_ALU_COMPARATOR_B1 enable_1/2_input_AND_5/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1289 enable_1/2_input_AND_5/OUT S0BAR_S1_DECODER enable_1/2_input_AND_5/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1290 VDD S0BAR_S1_DECODER enable_1/2_input_AND_6/OUT enable_1/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1291 enable_1/2_input_AND_6/a_4_n21# INPUT_ALU_B2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1292 OUTPUT_ALU_COMPARATOR_B2 enable_1/2_input_AND_6/OUT VDD enable_1/2_input_AND_6/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1293 enable_1/2_input_AND_6/OUT INPUT_ALU_B2 VDD enable_1/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 OUTPUT_ALU_COMPARATOR_B2 enable_1/2_input_AND_6/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1295 enable_1/2_input_AND_6/OUT S0BAR_S1_DECODER enable_1/2_input_AND_6/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1296 2_input_OR_0/OUT ADD_SUB_M GND Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1297 2_input_OR_0/a_n7_22# ADD_SUB_M VDD 2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1298 enable_2/enable 2_input_OR_0/OUT VDD 2_input_OR_0/w_30_15# CMOSP w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1299 enable_2/enable 2_input_OR_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=40 pd=26 as=0 ps=0
M1300 GND S0BAR_S1BAR_DECODER 2_input_OR_0/OUT Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 2_input_OR_0/OUT S0BAR_S1BAR_DECODER 2_input_OR_0/a_n7_22# 2_input_OR_0/w_n23_15# CMOSP w=4 l=2
+  ad=36 pd=26 as=0 ps=0
M1302 VDD enable_2/enable enable_2/2_input_AND_7/OUT enable_2/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1303 enable_2/2_input_AND_7/a_4_n21# INPUT_ALU_B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1304 OUTPUT_ALU_ADDER_B3 enable_2/2_input_AND_7/OUT VDD enable_2/2_input_AND_7/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1305 enable_2/2_input_AND_7/OUT INPUT_ALU_B3 VDD enable_2/2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1306 OUTPUT_ALU_ADDER_B3 enable_2/2_input_AND_7/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1307 enable_2/2_input_AND_7/OUT enable_2/enable enable_2/2_input_AND_7/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1308 VDD enable_2/enable enable_2/2_input_AND_0/OUT enable_2/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1309 enable_2/2_input_AND_0/a_4_n21# INPUT_ALU_A0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1310 OUTPUT_ALU_ADDER_A0 enable_2/2_input_AND_0/OUT VDD enable_2/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 enable_2/2_input_AND_0/OUT INPUT_ALU_A0 VDD enable_2/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 OUTPUT_ALU_ADDER_A0 enable_2/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1313 enable_2/2_input_AND_0/OUT enable_2/enable enable_2/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1314 VDD enable_2/enable enable_2/2_input_AND_1/OUT enable_2/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1315 enable_2/2_input_AND_1/a_4_n21# INPUT_ALU_A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1316 OUTPUT_ALU_ADDER_A1 enable_2/2_input_AND_1/OUT VDD enable_2/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1317 enable_2/2_input_AND_1/OUT INPUT_ALU_A1 VDD enable_2/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1318 OUTPUT_ALU_ADDER_A1 enable_2/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1319 enable_2/2_input_AND_1/OUT enable_2/enable enable_2/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1320 VDD enable_2/enable enable_2/2_input_AND_2/OUT enable_2/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1321 enable_2/2_input_AND_2/a_4_n21# INPUT_ALU_A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1322 OUTPUT_ALU_ADDER_A2 enable_2/2_input_AND_2/OUT VDD enable_2/2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1323 enable_2/2_input_AND_2/OUT INPUT_ALU_A2 VDD enable_2/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1324 OUTPUT_ALU_ADDER_A2 enable_2/2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1325 enable_2/2_input_AND_2/OUT enable_2/enable enable_2/2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1326 VDD enable_2/enable enable_2/2_input_AND_3/OUT enable_2/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1327 enable_2/2_input_AND_3/a_4_n21# INPUT_ALU_A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1328 OUTPUT_ALU_ADDER_A3 enable_2/2_input_AND_3/OUT VDD enable_2/2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1329 enable_2/2_input_AND_3/OUT INPUT_ALU_A3 VDD enable_2/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 OUTPUT_ALU_ADDER_A3 enable_2/2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1331 enable_2/2_input_AND_3/OUT enable_2/enable enable_2/2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1332 VDD enable_2/enable enable_2/2_input_AND_4/OUT enable_2/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1333 enable_2/2_input_AND_4/a_4_n21# INPUT_ALU_B0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1334 OUTPUT_ALU_ADDER_B0 enable_2/2_input_AND_4/OUT VDD enable_2/2_input_AND_4/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1335 enable_2/2_input_AND_4/OUT INPUT_ALU_B0 VDD enable_2/2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 OUTPUT_ALU_ADDER_B0 enable_2/2_input_AND_4/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1337 enable_2/2_input_AND_4/OUT enable_2/enable enable_2/2_input_AND_4/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1338 VDD enable_2/enable enable_2/2_input_AND_5/OUT enable_2/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1339 enable_2/2_input_AND_5/a_4_n21# INPUT_ALU_B1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1340 OUTPUT_ALU_ADDER_B1 enable_2/2_input_AND_5/OUT VDD enable_2/2_input_AND_5/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1341 enable_2/2_input_AND_5/OUT INPUT_ALU_B1 VDD enable_2/2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 OUTPUT_ALU_ADDER_B1 enable_2/2_input_AND_5/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1343 enable_2/2_input_AND_5/OUT enable_2/enable enable_2/2_input_AND_5/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1344 VDD enable_2/enable enable_2/2_input_AND_6/OUT enable_2/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1345 enable_2/2_input_AND_6/a_4_n21# INPUT_ALU_B2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1346 OUTPUT_ALU_ADDER_B2 enable_2/2_input_AND_6/OUT VDD enable_2/2_input_AND_6/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1347 enable_2/2_input_AND_6/OUT INPUT_ALU_B2 VDD enable_2/2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1348 OUTPUT_ALU_ADDER_B2 enable_2/2_input_AND_6/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1349 enable_2/2_input_AND_6/OUT enable_2/enable enable_2/2_input_AND_6/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1350 VDD COMPARATOR_OUT_A_EQUAL_B 2_input_AND_0/OUT 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1351 2_input_AND_0/a_4_n21# S0BAR_S1_DECODER GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1352 COMPARATOR_A_EQUAL_B_FINAL 2_input_AND_0/OUT VDD 2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1353 2_input_AND_0/OUT S0BAR_S1_DECODER VDD 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 COMPARATOR_A_EQUAL_B_FINAL 2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1355 2_input_AND_0/OUT COMPARATOR_OUT_A_EQUAL_B 2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1356 comparator_equal_0/B0_NOT OUTPUT_ALU_COMPARATOR_B0 VDD comparator_equal_0/q1a_NOT_3/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1357 comparator_equal_0/B0_NOT OUTPUT_ALU_COMPARATOR_B0 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1358 comparator_equal_0/q1a_NOT_4/out OUTPUT_ALU_COMPARATOR_A3 VDD comparator_equal_0/q1a_NOT_4/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1359 comparator_equal_0/q1a_NOT_4/out OUTPUT_ALU_COMPARATOR_A3 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1360 comparator_equal_0/A2NOT comparator_equal_0/q1a_NOT_5/in VDD comparator_equal_0/q1a_NOT_5/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1361 comparator_equal_0/A2NOT comparator_equal_0/q1a_NOT_5/in GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1362 comparator_equal_0/A0NOT OUTPUT_ALU_COMPARATOR_A0 VDD comparator_equal_0/q1a_NOT_6/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1363 comparator_equal_0/A0NOT OUTPUT_ALU_COMPARATOR_A0 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1364 comparator_equal_0/A1NOT OUTPUT_ALU_COMPARATOR_A1 VDD comparator_equal_0/q1a_NOT_7/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1365 comparator_equal_0/A1NOT OUTPUT_ALU_COMPARATOR_A1 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1366 VDD comparator_equal_0/A2B2 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=154 ps=86
M1367 comparator_equal_0/q1b_5_INPUT_AND_0/OUT OUTPUT_ALU_COMPARATOR_A0 VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1368 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A1B1 VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/q1b_5_INPUT_AND_0/OUT GND Gnd CMOSN w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1370 comparator_equal_0/q1b_5_INPUT_AND_0/a_n11_n43# comparator_equal_0/A3B3 GND Gnd CMOSN w=7 l=2
+  ad=56 pd=30 as=0 ps=0
M1371 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/q1b_5_INPUT_AND_0/OUT VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_50_10# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1372 comparator_equal_0/q1b_5_INPUT_AND_0/a_n1_n43# comparator_equal_0/A2B2 comparator_equal_0/q1b_5_INPUT_AND_0/a_n11_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1373 comparator_equal_0/q1b_5_INPUT_AND_0/OUT OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/q1b_5_INPUT_AND_0/a_17_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1374 comparator_equal_0/q1b_5_INPUT_AND_0/a_17_n43# comparator_equal_0/B0_NOT comparator_equal_0/q1b_5_INPUT_AND_0/a_8_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1375 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A3B3 VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 VDD comparator_equal_0/B0_NOT comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1377 comparator_equal_0/q1b_5_INPUT_AND_0/a_8_n43# comparator_equal_0/A1B1 comparator_equal_0/q1b_5_INPUT_AND_0/a_n1_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 VDD comparator_equal_0/A2B2 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=154 ps=86
M1379 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A0NOT VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A1B1 VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1b_5_INPUT_AND_1/OUT GND Gnd CMOSN w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1382 comparator_equal_0/q1b_5_INPUT_AND_1/a_n11_n43# comparator_equal_0/A3B3 GND Gnd CMOSN w=7 l=2
+  ad=56 pd=30 as=0 ps=0
M1383 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1b_5_INPUT_AND_1/OUT VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_50_10# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1384 comparator_equal_0/q1b_5_INPUT_AND_1/a_n1_n43# comparator_equal_0/A2B2 comparator_equal_0/q1b_5_INPUT_AND_1/a_n11_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1385 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A0NOT comparator_equal_0/q1b_5_INPUT_AND_1/a_17_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1386 comparator_equal_0/q1b_5_INPUT_AND_1/a_17_n43# OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/q1b_5_INPUT_AND_1/a_8_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1387 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A3B3 VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1388 VDD OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1389 comparator_equal_0/q1b_5_INPUT_AND_1/a_8_n43# comparator_equal_0/A1B1 comparator_equal_0/q1b_5_INPUT_AND_1/a_n1_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1390 COMPARATOR_OUT_A_GREATERTHAN_B comparator_equal_0/q1c_4_INPUT_OR_0/OUT VDD comparator_equal_0/q1c_4_INPUT_OR_0/w_41_n9# CMOSP w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1391 GND comparator_equal_0/A3_B3NOT comparator_equal_0/q1c_4_INPUT_OR_0/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=270 ps=114
M1392 comparator_equal_0/q1c_4_INPUT_OR_0/OUT comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/q1c_4_INPUT_OR_0/a_1_0# comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=90 pd=38 as=90 ps=38
M1393 comparator_equal_0/q1c_4_INPUT_OR_0/OUT comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1394 comparator_equal_0/q1c_4_INPUT_OR_0/OUT comparator_equal_0/A2_B2NOT_A3B3XNOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1395 comparator_equal_0/q1c_4_INPUT_OR_0/a_n18_0# comparator_equal_0/A3_B3NOT VDD comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1396 comparator_equal_0/q1c_4_INPUT_OR_0/a_1_0# comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/q1c_4_INPUT_OR_0/a_n9_0# comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1397 COMPARATOR_OUT_A_GREATERTHAN_B comparator_equal_0/q1c_4_INPUT_OR_0/OUT GND Gnd CMOSN w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1398 comparator_equal_0/q1c_4_INPUT_OR_0/a_n9_0# comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/q1c_4_INPUT_OR_0/a_n18_0# comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 GND comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/q1c_4_INPUT_OR_0/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1400 COMPARATOR_OUT_A_LESSTHAN_B comparator_equal_0/q1c_4_INPUT_OR_1/OUT VDD comparator_equal_0/q1c_4_INPUT_OR_1/w_41_n9# CMOSP w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1401 GND comparator_equal_0/A3NOT_B3 comparator_equal_0/q1c_4_INPUT_OR_1/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=270 ps=114
M1402 comparator_equal_0/q1c_4_INPUT_OR_1/OUT comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1c_4_INPUT_OR_1/a_1_0# comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=90 pd=38 as=90 ps=38
M1403 comparator_equal_0/q1c_4_INPUT_OR_1/OUT comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1404 comparator_equal_0/q1c_4_INPUT_OR_1/OUT comparator_equal_0/A2NOT_B2_A3B3XNOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 comparator_equal_0/q1c_4_INPUT_OR_1/a_n18_0# comparator_equal_0/A3NOT_B3 VDD comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1406 comparator_equal_0/q1c_4_INPUT_OR_1/a_1_0# comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1c_4_INPUT_OR_1/a_n9_0# comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1407 COMPARATOR_OUT_A_LESSTHAN_B comparator_equal_0/q1c_4_INPUT_OR_1/OUT GND Gnd CMOSN w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1408 comparator_equal_0/q1c_4_INPUT_OR_1/a_n9_0# comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/q1c_4_INPUT_OR_1/a_n18_0# comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 GND comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1c_4_INPUT_OR_1/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 comparator_equal_0/4_input_AND_0/a_n8_n45# comparator_equal_0/A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1411 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A2B2 VDD comparator_equal_0/4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=0 ps=0
M1412 COMPARATOR_OUT_A_EQUAL_B comparator_equal_0/4_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1413 VDD comparator_equal_0/A3B3 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1414 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A0B0 comparator_equal_0/4_input_AND_0/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1415 VDD comparator_equal_0/A1B1 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1416 COMPARATOR_OUT_A_EQUAL_B comparator_equal_0/4_input_AND_0/OUT VDD comparator_equal_0/4_input_AND_0/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1417 comparator_equal_0/4_input_AND_0/a_10_n45# comparator_equal_0/A1B1 comparator_equal_0/4_input_AND_0/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1418 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A0B0 VDD comparator_equal_0/4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 comparator_equal_0/4_input_AND_0/a_1_n45# comparator_equal_0/A2B2 comparator_equal_0/4_input_AND_0/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1420 comparator_equal_0/3_input_AND_0/OUT OUTPUT_ALU_COMPARATOR_A2 comparator_equal_0/3_input_AND_0/a_6_n34# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=24 ps=20
M1421 comparator_equal_0/3_input_AND_0/OUT OUTPUT_ALU_COMPARATOR_A2 VDD comparator_equal_0/3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=56 pd=44 as=0 ps=0
M1422 comparator_equal_0/3_input_AND_0/a_6_n34# comparator_equal_0/B2_NOT comparator_equal_0/3_input_AND_0/a_n3_n34# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=28 ps=22
M1423 VDD comparator_equal_0/B2_NOT comparator_equal_0/3_input_AND_0/OUT comparator_equal_0/3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 comparator_equal_0/3_input_AND_0/OUT comparator_equal_0/A3B3 VDD comparator_equal_0/3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1425 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/3_input_AND_0/OUT VDD comparator_equal_0/3_input_AND_0/w_34_3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1426 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/3_input_AND_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1427 comparator_equal_0/3_input_AND_0/a_n3_n34# comparator_equal_0/A3B3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 comparator_equal_0/4_input_AND_1/a_n8_n45# comparator_equal_0/A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1429 comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/A2B2 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=142 ps=96
M1430 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/4_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1431 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/A3B3 comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 comparator_equal_0/4_input_AND_1/OUT OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/4_input_AND_1/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1433 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/B1_NOT comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1434 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/4_input_AND_1/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1435 comparator_equal_0/4_input_AND_1/a_10_n45# comparator_equal_0/B1_NOT comparator_equal_0/4_input_AND_1/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1436 comparator_equal_0/4_input_AND_1/OUT OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1437 comparator_equal_0/4_input_AND_1/a_1_n45# comparator_equal_0/A2B2 comparator_equal_0/4_input_AND_1/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1438 VDD OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1439 comparator_equal_0/XNOR_1/OUT comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1440 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_B1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1441 VDD OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 comparator_equal_0/XNOR_1/OUT OUTPUT_ALU_COMPARATOR_B1 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1443 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_COMPARATOR_A1 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1444 comparator_equal_0/XNOR_1/OUT comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_A1 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1445 comparator_equal_0/XNOR_1/OUT OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1446 comparator_equal_0/A1B1 comparator_equal_0/XNOR_1/OUT VDD comparator_equal_0/XNOR_1/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1447 comparator_equal_0/A1B1 comparator_equal_0/XNOR_1/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1448 VDD OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1449 comparator_equal_0/XNOR_0/OUT comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1450 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_B0 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1451 VDD OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 comparator_equal_0/XNOR_0/OUT OUTPUT_ALU_COMPARATOR_B0 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1453 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_COMPARATOR_A0 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1454 comparator_equal_0/XNOR_0/OUT comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_A0 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1455 comparator_equal_0/XNOR_0/OUT OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1456 comparator_equal_0/A0B0 comparator_equal_0/XNOR_0/OUT VDD comparator_equal_0/XNOR_0/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1457 comparator_equal_0/A0B0 comparator_equal_0/XNOR_0/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1458 VDD OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/2_input_AND_0/OUT comparator_equal_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1459 comparator_equal_0/2_input_AND_0/a_4_n21# comparator_equal_0/B3_NOT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1460 comparator_equal_0/A3_B3NOT comparator_equal_0/2_input_AND_0/OUT VDD comparator_equal_0/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1461 comparator_equal_0/2_input_AND_0/OUT comparator_equal_0/B3_NOT VDD comparator_equal_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1462 comparator_equal_0/A3_B3NOT comparator_equal_0/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1463 comparator_equal_0/2_input_AND_0/OUT OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1464 comparator_equal_0/3_input_AND_1/OUT comparator_equal_0/A2NOT comparator_equal_0/3_input_AND_1/a_6_n34# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=24 ps=20
M1465 comparator_equal_0/3_input_AND_1/OUT comparator_equal_0/A2NOT VDD comparator_equal_0/3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=56 pd=44 as=0 ps=0
M1466 comparator_equal_0/3_input_AND_1/a_6_n34# OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/3_input_AND_1/a_n3_n34# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=28 ps=22
M1467 VDD OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/3_input_AND_1/OUT comparator_equal_0/3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 comparator_equal_0/3_input_AND_1/OUT comparator_equal_0/A3B3 VDD comparator_equal_0/3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1469 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/3_input_AND_1/OUT VDD comparator_equal_0/3_input_AND_1/w_34_3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1470 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/3_input_AND_1/OUT GND Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1471 comparator_equal_0/3_input_AND_1/a_n3_n34# comparator_equal_0/A3B3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 comparator_equal_0/4_input_AND_2/a_n8_n45# comparator_equal_0/A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1473 comparator_equal_0/4_input_AND_2/OUT comparator_equal_0/A2B2 VDD comparator_equal_0/4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=0 ps=0
M1474 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/4_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1475 VDD comparator_equal_0/A3B3 comparator_equal_0/4_input_AND_2/OUT comparator_equal_0/4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 comparator_equal_0/4_input_AND_2/OUT comparator_equal_0/A1NOT comparator_equal_0/4_input_AND_2/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1477 VDD OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/4_input_AND_2/OUT comparator_equal_0/4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1478 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/4_input_AND_2/OUT VDD comparator_equal_0/4_input_AND_2/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1479 comparator_equal_0/4_input_AND_2/a_10_n45# OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/4_input_AND_2/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1480 comparator_equal_0/4_input_AND_2/OUT comparator_equal_0/A1NOT VDD comparator_equal_0/4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1481 comparator_equal_0/4_input_AND_2/a_1_n45# comparator_equal_0/A2B2 comparator_equal_0/4_input_AND_2/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 VDD OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1483 comparator_equal_0/XNOR_2/OUT comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1484 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_B2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1485 VDD OUTPUT_ALU_COMPARATOR_A2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1486 comparator_equal_0/XNOR_2/OUT OUTPUT_ALU_COMPARATOR_B2 OUTPUT_ALU_COMPARATOR_A2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1487 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_COMPARATOR_A2 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1488 comparator_equal_0/XNOR_2/OUT comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_A2 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1489 comparator_equal_0/XNOR_2/OUT OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1490 comparator_equal_0/A2B2 comparator_equal_0/XNOR_2/OUT VDD comparator_equal_0/XNOR_2/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1491 comparator_equal_0/A2B2 comparator_equal_0/XNOR_2/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1492 VDD comparator_equal_0/q1a_NOT_4/out comparator_equal_0/2_input_AND_1/OUT comparator_equal_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1493 comparator_equal_0/2_input_AND_1/a_4_n21# OUTPUT_ALU_COMPARATOR_B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1494 comparator_equal_0/A3NOT_B3 comparator_equal_0/2_input_AND_1/OUT VDD comparator_equal_0/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1495 comparator_equal_0/2_input_AND_1/OUT OUTPUT_ALU_COMPARATOR_B3 VDD comparator_equal_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 comparator_equal_0/A3NOT_B3 comparator_equal_0/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1497 comparator_equal_0/2_input_AND_1/OUT comparator_equal_0/q1a_NOT_4/out comparator_equal_0/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1498 VDD OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1499 comparator_equal_0/XNOR_3/OUT comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1500 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_B3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1501 VDD OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1502 comparator_equal_0/XNOR_3/OUT OUTPUT_ALU_COMPARATOR_B3 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1503 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_COMPARATOR_A3 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1504 comparator_equal_0/XNOR_3/OUT comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_A3 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=0 ps=0
M1505 comparator_equal_0/XNOR_3/OUT OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1506 comparator_equal_0/A3B3 comparator_equal_0/XNOR_3/OUT VDD comparator_equal_0/XNOR_3/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1507 comparator_equal_0/A3B3 comparator_equal_0/XNOR_3/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1508 comparator_equal_0/B3_NOT OUTPUT_ALU_COMPARATOR_B3 VDD comparator_equal_0/q1a_NOT_0/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1509 comparator_equal_0/B3_NOT OUTPUT_ALU_COMPARATOR_B3 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1510 comparator_equal_0/B2_NOT OUTPUT_ALU_COMPARATOR_B2 VDD comparator_equal_0/q1a_NOT_1/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1511 comparator_equal_0/B2_NOT OUTPUT_ALU_COMPARATOR_B2 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1512 comparator_equal_0/B1_NOT OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/q1a_NOT_2/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1513 comparator_equal_0/B1_NOT OUTPUT_ALU_COMPARATOR_B1 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1514 VDD decoder_0/A0_BAR decoder_0/2_input_AND_0/OUT decoder_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1515 decoder_0/2_input_AND_0/a_4_n21# decoder_0/A1_BAR GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1516 S0BAR_S1BAR_DECODER decoder_0/2_input_AND_0/OUT VDD decoder_0/2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1517 decoder_0/2_input_AND_0/OUT decoder_0/A1_BAR VDD decoder_0/2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 S0BAR_S1BAR_DECODER decoder_0/2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1519 decoder_0/2_input_AND_0/OUT decoder_0/A0_BAR decoder_0/2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1520 VDD S0_DECODER decoder_0/2_input_AND_1/OUT decoder_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1521 decoder_0/2_input_AND_1/a_4_n21# decoder_0/A1_BAR GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1522 ADD_SUB_M decoder_0/2_input_AND_1/OUT VDD decoder_0/2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1523 decoder_0/2_input_AND_1/OUT decoder_0/A1_BAR VDD decoder_0/2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 ADD_SUB_M decoder_0/2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 decoder_0/2_input_AND_1/OUT S0_DECODER decoder_0/2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1526 VDD S1_DECODER decoder_0/2_input_AND_2/OUT decoder_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1527 decoder_0/2_input_AND_2/a_4_n21# decoder_0/A0_BAR GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1528 S0BAR_S1_DECODER decoder_0/2_input_AND_2/OUT VDD decoder_0/2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1529 decoder_0/2_input_AND_2/OUT decoder_0/A0_BAR VDD decoder_0/2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 S0BAR_S1_DECODER decoder_0/2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1531 decoder_0/2_input_AND_2/OUT S1_DECODER decoder_0/2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1532 VDD S1_DECODER decoder_0/2_input_AND_3/OUT decoder_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1533 decoder_0/2_input_AND_3/a_4_n21# S0_DECODER GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1534 S0_S1_DECODER decoder_0/2_input_AND_3/OUT VDD decoder_0/2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1535 decoder_0/2_input_AND_3/OUT S0_DECODER VDD decoder_0/2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 S0_S1_DECODER decoder_0/2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1537 decoder_0/2_input_AND_3/OUT S1_DECODER decoder_0/2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1538 decoder_0/A0_BAR S0_DECODER VDD decoder_0/q1a_NOT_0/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1539 decoder_0/A0_BAR S0_DECODER GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1540 decoder_0/A1_BAR S1_DECODER VDD decoder_0/q1a_NOT_1/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1541 decoder_0/A1_BAR S1_DECODER GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
C0 VDD adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.03fF
C1 adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_1/AXORB 0.07fF
C2 OUTPUT_ALU_ADDER_A0 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 0.32fF
C3 VDD comparator_equal_0/XNOR_0/w_181_105# 0.06fF
C4 VDD adder_subtractor_0/full_adder_3/AXORB 0.43fF
C5 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_3/AXORB 0.08fF
C6 VDD adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.06fF
C7 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_C1 0.09fF
C8 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/B0_XOR 0.09fF
C9 and_block_0/2_input_AND_2/OUT VDD 0.06fF
C10 S0BAR_S1_DECODER INPUT_ALU_A0 0.65fF
C11 adder_subtractor_0/B3_XOR adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.19fF
C12 and_block_0/2_input_AND_2/OUT AND_OUTPUT_A2B2 0.05fF
C13 VDD comparator_equal_0/A3_B3NOT 0.02fF
C14 ADD_SUB_M INPUT_ALU_A2 0.58fF
C15 enable_0/2_input_AND_1/OUT S0_S1_DECODER 0.12fF
C16 comparator_equal_0/XNOR_3/OUT comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C17 GND enable_0/2_input_AND_4/OUT 0.04fF
C18 OUTPUT_ALU_ADDER_A1 comparator_equal_0/A3NOT_B3 0.20fF
C19 comparator_equal_0/B2_NOT comparator_equal_0/3_input_AND_0/OUT 0.08fF
C20 adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# VDD 0.06fF
C21 VDD OUTPUT_ALU_COMPARATOR_B1 1.09fF
C22 VDD enable_1/2_input_AND_2/OUT 0.06fF
C23 comparator_equal_0/B2_NOT OUTPUT_ALU_COMPARATOR_A2 0.38fF
C24 INPUT_ALU_B0 INPUT_ALU_B2 0.64fF
C25 enable_2/2_input_AND_5/w_n12_9# enable_2/2_input_AND_5/OUT 0.03fF
C26 enable_1/2_input_AND_7/w_35_9# OUTPUT_ALU_COMPARATOR_B3 0.03fF
C27 ADD_SUB_M adder_subtractor_0/B3_XOR 0.18fF
C28 VDD adder_subtractor_0/q1d_2_INPUT_XOR_1/w_12_2# 0.03fF
C29 comparator_equal_0/A0B0 comparator_equal_0/A2B2 0.35fF
C30 comparator_equal_0/A3_B3NOT comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.09fF
C31 decoder_0/2_input_AND_3/OUT decoder_0/2_input_AND_3/w_35_9# 0.08fF
C32 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR VDD 0.03fF
C33 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_12_2# adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C34 VDD INPUT_ALU_A2 0.64fF
C35 OUTPUT_ALU_COMPARATOR_A2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C36 GND adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR 0.04fF
C37 adder_subtractor_0/B0_XOR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_53_n17# 0.04fF
C38 INPUT_ALU_B0 S0BAR_S1BAR_DECODER 0.11fF
C39 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/A2B2 0.19fF
C40 comparator_equal_0/4_input_AND_2/w_n22_4# comparator_equal_0/A2B2 0.07fF
C41 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_ADDER_A3 0.09fF
C42 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.09fF
C43 INPUT_ALU_B0 decoder_0/2_input_AND_1/OUT 0.13fF
C44 S0BAR_S1_DECODER 2_input_AND_0/w_n12_9# 0.07fF
C45 S0_S1_DECODER INPUT_ALU_B2 0.75fF
C46 adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# adder_subtractor_0/B0_XOR 0.07fF
C47 enable_0/2_input_AND_7/w_n12_9# INPUT_ALU_B3 0.07fF
C48 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_53_n17# ADDER_SUB_CFINAL 0.04fF
C49 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_12_2# adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR 0.03fF
C50 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_n34_1# adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.03fF
C51 VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_50_10# 0.06fF
C52 VDD adder_subtractor_0/B3_XOR 1.22fF
C53 VDD adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.06fF
C54 and_block_0/2_input_AND_1/OUT VDD 0.06fF
C55 OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/4_input_AND_2/OUT 0.09fF
C56 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_53_n17# 0.09fF
C57 ADD_SUB_M INPUT_ALU_A0 0.30fF
C58 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_A1 0.19fF
C59 enable_2/enable enable_2/2_input_AND_0/w_n12_9# 0.07fF
C60 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C61 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C62 GND enable_2/enable 4.24fF
C63 adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.12fF
C64 S0BAR_S1_DECODER INPUT_ALU_B3 0.57fF
C65 OUTPUT_ALU_ADDER_A2 enable_2/2_input_AND_2/w_35_9# 0.03fF
C66 ADDER_SUB_S1 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR 0.19fF
C67 OUTPUT_ALU_COMPARATOR_A1 OUTPUT_ALU_COMPARATOR_B2 0.18fF
C68 GND enable_0/2_input_AND_3/OUT 0.04fF
C69 INPUT_ALU_A3 decoder_0/2_input_AND_0/OUT 0.37fF
C70 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# OUTPUT_ALU_ADDER_B1 0.09fF
C71 adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# VDD 0.03fF
C72 GND adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C73 INPUT_ALU_A3 INPUT_ALU_B2 0.72fF
C74 INPUT_ALU_B0 INPUT_ALU_B1 0.72fF
C75 VDD enable_0/2_input_AND_6/w_35_9# 0.03fF
C76 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR GND 0.08fF
C77 VDD INPUT_ALU_A0 0.64fF
C78 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT ADDER_SUB_C1 0.05fF
C79 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/A3B3 0.08fF
C80 comparator_equal_0/A1B1 comparator_equal_0/A2B2 4.95fF
C81 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/A3B3 0.08fF
C82 VDD enable_2/2_input_AND_6/w_n12_9# 0.07fF
C83 OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/q1a_NOT_2/w_n12_4# 0.10fF
C84 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/B1_NOT 0.37fF
C85 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_1/w_n34_1# 0.08fF
C86 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_B0 0.03fF
C87 VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# 0.15fF
C88 GND adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.04fF
C89 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/A3B3 4.76fF
C90 VDD decoder_0/q1a_NOT_0/w_n12_4# 0.08fF
C91 S0_S1_DECODER INPUT_ALU_B1 0.70fF
C92 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/4_input_AND_1/a_1_n45# 0.01fF
C93 adder_subtractor_0/full_adder_1/2_input_OR_0/A adder_subtractor_0/full_adder_1/2_input_AND_1/w_35_9# 0.03fF
C94 adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# adder_subtractor_0/B1_XOR 0.07fF
C95 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_C2 0.09fF
C96 GND comparator_equal_0/A2_B2NOT_A3B3XNOR 0.10fF
C97 VDD comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.32fF
C98 VDD adder_subtractor_0/full_adder_1/2_input_OR_0/OUT 0.02fF
C99 VDD adder_subtractor_0/full_adder_3/2_input_OR_0/B 0.12fF
C100 ADD_SUB_M decoder_0/2_input_AND_1/w_35_9# 0.03fF
C101 OUTPUT_ALU_ADDER_A3 OUTPUT_ALU_ADDER_B1 0.30fF
C102 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# comparator_equal_0/A1B1 0.07fF
C103 adder_subtractor_0/B1_XOR OUTPUT_ALU_ADDER_B1 0.22fF
C104 and_block_0/2_input_AND_0/OUT VDD 0.06fF
C105 ADD_SUB_M INPUT_ALU_B3 0.60fF
C106 comparator_equal_0/B1_NOT comparator_equal_0/A3B3 0.08fF
C107 VDD adder_subtractor_0/q1d_2_INPUT_XOR_1/w_n34_1# 0.03fF
C108 ADDER_SUB_S2 ADDER_SUB_C2 0.15fF
C109 adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.05fF
C110 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR ADD_SUB_M 0.51fF
C111 comparator_equal_0/4_input_AND_0/w_40_5# COMPARATOR_OUT_A_EQUAL_B 0.03fF
C112 and_block_0/2_input_AND_1/OUT AND_OUTPUT_A1B1 0.05fF
C113 INPUT_ALU_B2 OUTPUT_ALU_COMPARATOR_B1 0.04fF
C114 INPUT_ALU_A1 decoder_0/2_input_AND_2/w_35_9# 0.01fF
C115 GND comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.63fF
C116 GND comparator_equal_0/A1NOT 0.13fF
C117 VDD 2_input_AND_0/w_n12_9# 0.06fF
C118 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C119 comparator_equal_0/A1B1 comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.08fF
C120 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/A0NOT 1.29fF
C121 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/A0NOT 0.04fF
C122 GND adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR 0.04fF
C123 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_n34_1# 0.03fF
C124 INPUT_ALU_A3 decoder_0/A0_BAR 0.02fF
C125 VDD enable_0/2_input_AND_5/w_35_9# 0.03fF
C126 INPUT_ALU_A2 INPUT_ALU_B2 0.86fF
C127 INPUT_ALU_A3 INPUT_ALU_B1 0.68fF
C128 enable_2/2_input_AND_4/w_n12_9# enable_2/2_input_AND_4/OUT 0.03fF
C129 enable_1/2_input_AND_1/w_35_9# OUTPUT_ALU_COMPARATOR_A1 0.13fF
C130 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_12_2# adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR 0.03fF
C131 VDD 2_input_AND_0/w_35_9# 0.03fF
C132 VDD decoder_0/2_input_AND_1/w_35_9# 0.03fF
C133 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_12_2# ADDER_SUB_C3 0.08fF
C134 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR VDD 0.03fF
C135 VDD INPUT_ALU_B3 0.23fF
C136 VDD comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C137 VDD enable_2/2_input_AND_5/w_n12_9# 0.06fF
C138 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C139 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_n34_1# adder_subtractor_0/B1_XOR 0.08fF
C140 VDD comparator_equal_0/q1a_NOT_1/w_n12_4# 0.07fF
C141 GND adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.04fF
C142 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/A2NOT 0.39fF
C143 VDD comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C144 decoder_0/2_input_AND_2/OUT S1_DECODER 0.12fF
C145 enable_2/enable enable_2/2_input_AND_7/w_n12_9# 0.07fF
C146 S0_S1_DECODER INPUT_ALU_B0 0.72fF
C147 enable_1/2_input_AND_5/OUT OUTPUT_ALU_COMPARATOR_B1 0.05fF
C148 adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_0/2_input_OR_0/A 0.07fF
C149 OUTPUT_ALU_ADDER_B3 adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR 0.03fF
C150 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/q1a_NOT_2/w_n12_4# 0.05fF
C151 GND S1_DECODER 0.55fF
C152 VDD comparator_equal_0/q1a_NOT_4/out 0.46fF
C153 enable_0/2_input_AND_7/w_35_9# OUTPUT_ALU_ANDBLOCK_B3 0.03fF
C154 enable_0/2_input_AND_6/w_n12_9# enable_0/2_input_AND_6/OUT 0.03fF
C155 comparator_equal_0/B0_NOT OUTPUT_ALU_COMPARATOR_B0 0.04fF
C156 enable_0/2_input_AND_0/w_n12_9# S0_S1_DECODER 0.07fF
C157 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/B0_NOT 0.84fF
C158 enable_1/2_input_AND_3/w_35_9# OUTPUT_ALU_COMPARATOR_A3 0.13fF
C159 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C3 0.03fF
C160 ADDER_SUB_S3 adder_subtractor_0/full_adder_3/AXORB 0.18fF
C161 adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_OR_0/OUT 0.20fF
C162 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_53_n17# ADDER_SUB_S1 0.04fF
C163 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_1/AXORB 0.24fF
C164 GND decoder_0/2_input_AND_2/OUT 0.04fF
C165 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C166 INPUT_ALU_A0 INPUT_ALU_B2 0.56fF
C167 enable_2/2_input_AND_6/w_n12_9# INPUT_ALU_B2 0.07fF
C168 OUTPUT_ALU_ADDER_A1 enable_2/2_input_AND_1/w_35_9# 0.08fF
C169 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C170 S0BAR_S1_DECODER OUTPUT_ALU_COMPARATOR_A1 0.30fF
C171 INPUT_ALU_A2 decoder_0/A0_BAR 0.27fF
C172 comparator_equal_0/A2B2 comparator_equal_0/XNOR_2/w_181_105# 0.06fF
C173 INPUT_ALU_A3 INPUT_ALU_B0 0.65fF
C174 INPUT_ALU_A2 INPUT_ALU_B1 0.81fF
C175 VDD enable_0/2_input_AND_4/w_35_9# 0.03fF
C176 VDD enable_0/2_input_AND_1/w_35_9# 0.03fF
C177 VDD comparator_equal_0/4_input_AND_0/OUT 0.21fF
C178 VDD enable_2/2_input_AND_4/w_n12_9# 0.06fF
C179 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C180 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_12_2# ADD_SUB_M 0.08fF
C181 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# comparator_equal_0/A2NOT_B2_A3B3XNOR 0.10fF
C182 GND adder_subtractor_0/full_adder_3/2_input_OR_0/OUT 0.15fF
C183 decoder_0/2_input_AND_3/OUT S1_DECODER 0.12fF
C184 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C185 S0_S1_DECODER INPUT_ALU_A3 0.74fF
C186 OUTPUT_ALU_ANDBLOCK_A3 VDD 1.03fF
C187 adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_1/2_input_OR_0/B 0.07fF
C188 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.06fF
C189 adder_subtractor_0/full_adder_2/2_input_AND_1/w_35_9# adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.08fF
C190 ADDER_SUB_C2 adder_subtractor_0/full_adder_2/AXORB 0.93fF
C191 adder_subtractor_0/full_adder_0/AXORB adder_subtractor_0/full_adder_0/2_input_AND_1/OUT 0.12fF
C192 AND_OUTPUT_A2B2 OUTPUT_ALU_ANDBLOCK_A3 0.37fF
C193 comparator_equal_0/q1a_NOT_6/w_n12_4# comparator_equal_0/A0NOT 0.09fF
C194 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_12_2# VDD 0.03fF
C195 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_A2 0.08fF
C196 adder_subtractor_0/full_adder_3/2_input_OR_0/w_30_15# ADDER_SUB_C4 0.03fF
C197 OUTPUT_ALU_COMPARATOR_B0 OUTPUT_ALU_COMPARATOR_B3 0.54fF
C198 GND decoder_0/2_input_AND_3/OUT 0.04fF
C199 VDD comparator_equal_0/XNOR_1/w_181_105# 0.06fF
C200 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_B3 0.19fF
C201 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_2/AXORB 0.04fF
C202 INPUT_ALU_A0 INPUT_ALU_B1 0.52fF
C203 VDD comparator_equal_0/A2NOT_B2_A3B3XNOR 0.31fF
C204 GND comparator_equal_0/B2_NOT 0.12fF
C205 INPUT_ALU_B3 INPUT_ALU_B2 1.05fF
C206 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C207 GND adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR 0.27fF
C208 OUTPUT_ALU_COMPARATOR_B2 OUTPUT_ALU_COMPARATOR_B3 0.44fF
C209 and_block_0/2_input_AND_0/OUT AND_OUTPUT_A0B0 0.05fF
C210 INPUT_ALU_A2 INPUT_ALU_B0 0.80fF
C211 enable_2/2_input_AND_3/w_n12_9# enable_2/2_input_AND_3/OUT 0.03fF
C212 VDD adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.06fF
C213 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_12_2# OUTPUT_ALU_ADDER_A3 0.08fF
C214 VDD enable_2/2_input_AND_3/w_n12_9# 0.06fF
C215 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_12_2# VDD 0.03fF
C216 decoder_0/A0_BAR decoder_0/q1a_NOT_0/w_n12_4# 0.04fF
C217 GND comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.23fF
C218 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C219 decoder_0/2_input_AND_1/OUT decoder_0/2_input_AND_1/w_35_9# 0.08fF
C220 enable_0/2_input_AND_1/OUT enable_0/2_input_AND_1/w_35_9# 0.08fF
C221 decoder_0/q1a_NOT_1/w_n12_4# decoder_0/A1_BAR 0.04fF
C222 S0BAR_S1_DECODER enable_1/2_input_AND_6/w_n12_9# 0.07fF
C223 GND ADDER_SUB_S1 0.05fF
C224 adder_subtractor_0/B3_XOR adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# 0.03fF
C225 VDD OUTPUT_ALU_COMPARATOR_A1 1.67fF
C226 OUTPUT_ALU_ADDER_A0 comparator_equal_0/A3NOT_B3 0.32fF
C227 S0_S1_DECODER INPUT_ALU_A2 0.70fF
C228 VDD enable_0/2_input_AND_0/OUT 0.06fF
C229 VDD comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C230 OUTPUT_ALU_ANDBLOCK_A2 VDD 0.89fF
C231 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_2/w_n34_1# 0.08fF
C232 VDD adder_subtractor_0/full_adder_3/2_input_AND_1/w_35_9# 0.03fF
C233 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_1/AXORB 0.08fF
C234 VDD ADDER_SUB_C1 0.15fF
C235 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_A3 0.20fF
C236 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# comparator_equal_0/XNOR_3/OUT 0.03fF
C237 ADDER_SUB_C4 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_n34_1# 0.08fF
C238 OUTPUT_ALU_ADDER_A2 adder_subtractor_0/full_adder_2/AXORB 0.15fF
C239 VDD comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# 0.11fF
C240 enable_0/2_input_AND_5/w_n12_9# enable_0/2_input_AND_5/OUT 0.03fF
C241 VDD comparator_equal_0/2_input_AND_0/w_n12_9# 0.06fF
C242 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_n34_1# OUTPUT_ALU_ADDER_A0 0.08fF
C243 enable_1/2_input_AND_0/w_n12_9# INPUT_ALU_A0 0.07fF
C244 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR 0.09fF
C245 INPUT_ALU_A0 INPUT_ALU_B0 0.51fF
C246 comparator_equal_0/2_input_AND_0/w_35_9# comparator_equal_0/2_input_AND_0/OUT 0.08fF
C247 comparator_equal_0/B3_NOT comparator_equal_0/2_input_AND_0/w_n12_9# 0.07fF
C248 comparator_equal_0/3_input_AND_0/w_34_3# comparator_equal_0/3_input_AND_0/OUT 0.06fF
C249 GND enable_0/2_input_AND_7/OUT 0.04fF
C250 VDD comparator_equal_0/A3B3 2.00fF
C251 VDD enable_0/2_input_AND_2/OUT 0.06fF
C252 INPUT_ALU_B3 INPUT_ALU_B1 1.02fF
C253 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_COMPARATOR_A2 0.03fF
C254 enable_2/2_input_AND_5/w_n12_9# INPUT_ALU_B1 0.07fF
C255 VDD adder_subtractor_0/q1d_2_INPUT_XOR_2/w_n34_1# 0.03fF
C256 enable_1/2_input_AND_7/OUT OUTPUT_ALU_COMPARATOR_B3 0.05fF
C257 ADD_SUB_M OUTPUT_ALU_ADDER_A1 0.31fF
C258 INPUT_ALU_A2 INPUT_ALU_A3 1.17fF
C259 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.10fF
C260 comparator_equal_0/q1b_5_INPUT_AND_1/w_50_10# comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.04fF
C261 OUTPUT_ALU_ADDER_A2 OUTPUT_ALU_ADDER_B2 0.39fF
C262 VDD adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.06fF
C263 enable_0/2_input_AND_0/w_n12_9# INPUT_ALU_A0 0.07fF
C264 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# 0.09fF
C265 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C266 OUTPUT_ALU_COMPARATOR_A2 comparator_equal_0/XNOR_2/OUT 0.18fF
C267 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C268 VDD enable_2/2_input_AND_2/w_n12_9# 0.06fF
C269 GND OUTPUT_ALU_ADDER_B3 0.91fF
C270 S0_S1_DECODER INPUT_ALU_A0 0.59fF
C271 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_A3 0.08fF
C272 adder_subtractor_0/B0_XOR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C273 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_ADDER_A1 0.09fF
C274 OUTPUT_ALU_COMPARATOR_A0 INPUT_ALU_A1 0.03fF
C275 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/A2B2 0.29fF
C276 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/A3B3 1.07fF
C277 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/3_input_AND_1/w_34_3# 0.03fF
C278 comparator_equal_0/q1c_4_INPUT_OR_0/w_41_n9# comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.10fF
C279 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A1 0.03fF
C280 S0BAR_S1_DECODER enable_1/2_input_AND_5/w_n12_9# 0.07fF
C281 comparator_equal_0/XNOR_2/OUT comparator_equal_0/XNOR_2/w_181_105# 0.13fF
C282 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_53_n17# 0.09fF
C283 VDD OUTPUT_ALU_ADDER_A1 1.38fF
C284 comparator_equal_0/A2B2 comparator_equal_0/A1NOT 0.08fF
C285 comparator_equal_0/A3B3 comparator_equal_0/4_input_AND_2/OUT 0.15fF
C286 OUTPUT_ALU_ANDBLOCK_A1 VDD 0.95fF
C287 VDD adder_subtractor_0/full_adder_3/2_input_AND_0/w_35_9# 0.03fF
C288 2_input_AND_0/w_n12_9# COMPARATOR_OUT_A_EQUAL_B 0.07fF
C289 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/OUT 0.15fF
C290 adder_subtractor_0/full_adder_2/2_input_AND_0/w_35_9# adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.08fF
C291 OUTPUT_ALU_ADDER_A2 adder_subtractor_0/B2_XOR 1.32fF
C292 OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT 0.12fF
C293 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/OUT 0.18fF
C294 adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/AXORB 0.18fF
C295 GND comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 0.06fF
C296 VDD comparator_equal_0/A0NOT 0.10fF
C297 VDD enable_1/2_input_AND_6/w_n12_9# 0.07fF
C298 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_ADDER_B0 0.09fF
C299 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR OUTPUT_ALU_ADDER_B1 0.08fF
C300 INPUT_ALU_A0 INPUT_ALU_A3 0.89fF
C301 comparator_equal_0/q1a_NOT_4/out comparator_equal_0/2_input_AND_1/OUT 0.12fF
C302 adder_subtractor_0/B1_XOR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_53_n17# 0.04fF
C303 INPUT_ALU_B0 decoder_0/2_input_AND_1/w_35_9# 0.02fF
C304 GND COMPARATOR_OUT_A_LESSTHAN_B 0.04fF
C305 VDD comparator_equal_0/A2NOT 0.10fF
C306 INPUT_ALU_B3 INPUT_ALU_B0 0.91fF
C307 ADD_SUB_M 2_input_OR_0/w_n23_15# 0.07fF
C308 adder_subtractor_0/full_adder_1/2_input_OR_0/w_30_15# ADDER_SUB_C2 0.03fF
C309 comparator_equal_0/A0B0 OUTPUT_ALU_COMPARATOR_B2 0.32fF
C310 enable_2/2_input_AND_2/w_n12_9# enable_2/2_input_AND_2/OUT 0.03fF
C311 VDD adder_subtractor_0/full_adder_2/2_input_OR_0/OUT 0.02fF
C312 VDD OUTPUT_ALU_ANDBLOCK_B2 0.91fF
C313 GND adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR 0.04fF
C314 GND ADDER_SUB_C3 0.80fF
C315 GND adder_subtractor_0/full_adder_1/AXORB 0.33fF
C316 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR OUTPUT_ALU_COMPARATOR_B2 0.42fF
C317 S0BAR_S1_DECODER enable_1/2_input_AND_4/w_n12_9# 0.07fF
C318 S0_S1_DECODER INPUT_ALU_B3 0.55fF
C319 VDD comparator_equal_0/B0_NOT 0.10fF
C320 GND comparator_equal_0/2_input_AND_0/OUT 0.04fF
C321 VDD 2_input_OR_0/w_n23_15# 0.03fF
C322 VDD adder_subtractor_0/full_adder_3/2_input_OR_0/w_30_15# 0.03fF
C323 VDD adder_subtractor_0/full_adder_1/2_input_OR_0/A 0.18fF
C324 OUTPUT_ALU_ADDER_A1 OUTPUT_ALU_ADDER_B0 0.22fF
C325 OUTPUT_ALU_ANDBLOCK_A0 VDD 0.93fF
C326 ADDER_SUB_S0 ADD_SUB_M 0.15fF
C327 adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_AND_0/OUT 0.05fF
C328 comparator_equal_0/4_input_AND_0/w_40_5# comparator_equal_0/4_input_AND_0/OUT 0.07fF
C329 OUTPUT_ALU_ANDBLOCK_A1 enable_0/2_input_AND_1/OUT 0.05fF
C330 adder_subtractor_0/full_adder_3/2_input_OR_0/A adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.05fF
C331 GND comparator_equal_0/A2B2 1.52fF
C332 VDD 2_input_OR_0/w_30_15# 0.03fF
C333 enable_0/2_input_AND_4/w_n12_9# enable_0/2_input_AND_4/OUT 0.03fF
C334 VDD enable_0/2_input_AND_2/w_35_9# 0.03fF
C335 VDD enable_1/2_input_AND_5/w_n12_9# 0.06fF
C336 comparator_equal_0/A1B1 OUTPUT_ALU_COMPARATOR_B0 1.08fF
C337 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/A1B1 0.08fF
C338 INPUT_ALU_A0 INPUT_ALU_A2 0.76fF
C339 S0BAR_S1_DECODER OUTPUT_ALU_COMPARATOR_A3 0.29fF
C340 comparator_equal_0/4_input_AND_0/OUT COMPARATOR_OUT_A_EQUAL_B 0.04fF
C341 comparator_equal_0/q1a_NOT_5/in comparator_equal_0/A3B3 1.07fF
C342 INPUT_ALU_B3 INPUT_ALU_A3 0.65fF
C343 enable_2/2_input_AND_4/w_n12_9# INPUT_ALU_B0 0.07fF
C344 INPUT_ALU_A1 S0_DECODER 0.07fF
C345 VDD 2_input_AND_0/OUT 0.06fF
C346 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_12_2# ADDER_SUB_C1 0.08fF
C347 comparator_equal_0/A1B1 OUTPUT_ALU_COMPARATOR_B2 0.84fF
C348 VDD comparator_equal_0/3_input_AND_0/w_n19_2# 0.06fF
C349 VDD enable_1/2_input_AND_2/w_35_9# 0.03fF
C350 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR 0.03fF
C351 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_12_2# OUTPUT_ALU_ADDER_B2 0.08fF
C352 VDD OUTPUT_ALU_ANDBLOCK_B1 0.87fF
C353 INPUT_ALU_A2 decoder_0/q1a_NOT_0/w_n12_4# 0.03fF
C354 OUTPUT_ALU_ANDBLOCK_A3 INPUT_ALU_B0 0.04fF
C355 VDD comparator_equal_0/XNOR_3/w_181_105# 0.06fF
C356 enable_1/2_input_AND_6/w_n12_9# enable_1/2_input_AND_6/OUT 0.03fF
C357 GND OUTPUT_ALU_ADDER_A3 0.73fF
C358 GND adder_subtractor_0/B1_XOR 0.73fF
C359 comparator_equal_0/3_input_AND_1/w_n19_2# comparator_equal_0/3_input_AND_1/OUT 0.06fF
C360 VDD adder_subtractor_0/q1d_2_INPUT_XOR_4/w_n34_1# 0.03fF
C361 OUTPUT_ALU_ADDER_A1 enable_2/2_input_AND_1/OUT 0.05fF
C362 S0BAR_S1_DECODER enable_1/2_input_AND_3/w_n12_9# 0.07fF
C363 S1_DECODER decoder_0/2_input_AND_2/w_n12_9# 0.07fF
C364 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/3_input_AND_0/w_34_3# 0.03fF
C365 GND comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.06fF
C366 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.03fF
C367 VDD OUTPUT_ALU_COMPARATOR_B3 3.38fF
C368 decoder_0/2_input_AND_2/OUT decoder_0/2_input_AND_2/w_n12_9# 0.03fF
C369 enable_1/2_input_AND_6/w_n12_9# INPUT_ALU_B2 0.07fF
C370 VDD adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR 0.03fF
C371 S0BAR_S1_DECODER INPUT_ALU_A1 0.75fF
C372 adder_subtractor_0/full_adder_2/2_input_OR_0/A adder_subtractor_0/full_adder_2/2_input_OR_0/B 0.45fF
C373 adder_subtractor_0/full_adder_2/2_input_OR_0/w_30_15# adder_subtractor_0/full_adder_2/2_input_OR_0/OUT 0.06fF
C374 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C1 0.03fF
C375 ADDER_SUB_S1 adder_subtractor_0/full_adder_1/AXORB 0.18fF
C376 adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_OR_0/OUT 0.20fF
C377 GND comparator_equal_0/3_input_AND_1/OUT 0.09fF
C378 enable_0/2_input_AND_0/OUT enable_0/2_input_AND_0/w_35_9# 0.08fF
C379 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_1/OUT 0.04fF
C380 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C381 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C382 comparator_equal_0/B3_NOT OUTPUT_ALU_COMPARATOR_B3 0.04fF
C383 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_S3 0.03fF
C384 AND_OUTPUT_A0B0 OUTPUT_ALU_ANDBLOCK_A1 0.30fF
C385 VDD enable_1/2_input_AND_4/w_n12_9# 0.06fF
C386 comparator_equal_0/q1a_NOT_7/w_n12_4# comparator_equal_0/A1NOT 0.04fF
C387 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR OUTPUT_ALU_COMPARATOR_B3 0.59fF
C388 comparator_equal_0/q1a_NOT_5/in comparator_equal_0/A2NOT 0.04fF
C389 OUTPUT_ALU_ADDER_B3 enable_2/2_input_AND_7/w_35_9# 0.03fF
C390 INPUT_ALU_B3 INPUT_ALU_A2 0.79fF
C391 comparator_equal_0/4_input_AND_1/w_40_5# comparator_equal_0/4_input_AND_1/OUT 0.07fF
C392 comparator_equal_0/4_input_AND_1/w_n22_4# comparator_equal_0/q1a_NOT_2/vdd 0.05fF
C393 GND comparator_equal_0/4_input_AND_1/OUT 0.11fF
C394 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C395 VDD OUTPUT_ALU_ANDBLOCK_B0 3.56fF
C396 GND adder_subtractor_0/full_adder_3/2_input_OR_0/A 0.44fF
C397 GND adder_subtractor_0/full_adder_1/2_input_OR_0/B 0.16fF
C398 OUTPUT_ALU_COMPARATOR_A0 enable_1/2_input_AND_0/OUT 0.05fF
C399 VDD OUTPUT_ALU_COMPARATOR_A3 1.13fF
C400 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.08fF
C401 and_block_0/2_input_AND_3/w_n12_9# VDD 0.06fF
C402 comparator_equal_0/4_input_AND_0/w_n22_4# comparator_equal_0/A2B2 0.07fF
C403 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C404 VDD comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C405 OUTPUT_ALU_ADDER_B1 enable_2/2_input_AND_5/OUT 0.05fF
C406 enable_0/2_input_AND_0/OUT enable_0/2_input_AND_0/w_n12_9# 0.03fF
C407 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_A2 0.21fF
C408 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/B3_NOT 0.57fF
C409 adder_subtractor_0/full_adder_0/2_input_AND_1/w_35_9# adder_subtractor_0/full_adder_0/2_input_AND_1/OUT 0.08fF
C410 ADD_SUB_M adder_subtractor_0/full_adder_0/AXORB 0.93fF
C411 ADD_SUB_M INPUT_ALU_A1 0.53fF
C412 GND COMPARATOR_A_EQUAL_B_FINAL 0.05fF
C413 2_input_OR_0/w_n23_15# S0BAR_S1BAR_DECODER 0.07fF
C414 VDD enable_0/2_input_AND_2/w_n12_9# 0.06fF
C415 adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_2/AXORB 0.07fF
C416 enable_0/2_input_AND_0/OUT S0_S1_DECODER 0.12fF
C417 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.78fF
C418 decoder_0/A1_BAR S1_DECODER 0.04fF
C419 OUTPUT_ALU_COMPARATOR_B2 OUTPUT_ALU_COMPARATOR_A2 0.76fF
C420 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.42fF
C421 VDD comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C422 decoder_0/2_input_AND_2/OUT decoder_0/2_input_AND_2/w_35_9# 0.08fF
C423 INPUT_ALU_B3 INPUT_ALU_A0 0.51fF
C424 VDD enable_1/2_input_AND_3/w_n12_9# 0.06fF
C425 VDD comparator_equal_0/q1c_4_INPUT_OR_1/w_41_n9# 0.20fF
C426 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_0/OUT 0.04fF
C427 GND ADDER_SUB_S2 0.05fF
C428 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR GND 0.04fF
C429 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_12_2# VDD 0.03fF
C430 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_n34_1# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C431 enable_2/2_input_AND_3/w_n12_9# INPUT_ALU_A3 0.07fF
C432 enable_1/2_input_AND_1/w_35_9# enable_1/2_input_AND_1/OUT 0.08fF
C433 VDD ADDER_SUB_C2 0.15fF
C434 adder_subtractor_0/full_adder_0/AXORB VDD 0.43fF
C435 VDD INPUT_ALU_A1 0.38fF
C436 GND decoder_0/A1_BAR 0.20fF
C437 enable_0/2_input_AND_2/OUT S0_S1_DECODER 0.12fF
C438 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C439 VDD OUTPUT_ALU_ANDBLOCK_B3 0.83fF
C440 2_input_OR_0/w_n23_15# INPUT_ALU_B1 0.02fF
C441 enable_1/2_input_AND_5/w_n12_9# enable_1/2_input_AND_5/OUT 0.03fF
C442 GND adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.18fF
C443 VDD adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# 0.06fF
C444 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_12_2# adder_subtractor_0/B0_XOR 0.08fF
C445 and_block_0/2_input_AND_2/w_n12_9# VDD 0.06fF
C446 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/A2B2 0.25fF
C447 VDD comparator_equal_0/XNOR_0/OUT 0.17fF
C448 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_3/AXORB 0.04fF
C449 2_input_OR_0/w_30_15# INPUT_ALU_B1 0.02fF
C450 comparator_equal_0/q1a_NOT_3/w_n12_4# OUTPUT_ALU_COMPARATOR_B0 0.09fF
C451 VDD enable_0/2_input_AND_3/w_35_9# 0.03fF
C452 OUTPUT_ALU_ADDER_A3 OUTPUT_ALU_ADDER_B3 0.36fF
C453 ADD_SUB_M OUTPUT_ALU_ADDER_A2 0.49fF
C454 OUTPUT_ALU_ADDER_A0 ADD_SUB_M 0.52fF
C455 comparator_equal_0/q1a_NOT_5/in OUTPUT_ALU_COMPARATOR_B3 0.28fF
C456 adder_subtractor_0/B0_XOR adder_subtractor_0/full_adder_0/AXORB 0.15fF
C457 enable_1/2_input_AND_5/w_n12_9# INPUT_ALU_B1 0.07fF
C458 adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.03fF
C459 VDD comparator_equal_0/A0B0 0.42fF
C460 VDD adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C461 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR VDD 0.03fF
C462 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_52_34# adder_subtractor_0/full_adder_3/AXORB 0.03fF
C463 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C464 VDD comparator_equal_0/4_input_AND_2/w_n22_4# 0.05fF
C465 VDD comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.07fF
C466 OUTPUT_ALU_ANDBLOCK_A0 enable_0/2_input_AND_0/w_35_9# 0.12fF
C467 S0BAR_S1_DECODER enable_1/2_input_AND_1/OUT 0.12fF
C468 ADDER_SUB_S2 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR 0.19fF
C469 GND adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C470 OUTPUT_ALU_COMPARATOR_A1 OUTPUT_ALU_COMPARATOR_B1 0.52fF
C471 OUTPUT_ALU_ADDER_A1 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.19fF
C472 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# comparator_equal_0/A3_B3NOT 0.12fF
C473 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_n34_1# adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.03fF
C474 VDD OUTPUT_ALU_ADDER_A2 1.03fF
C475 OUTPUT_ALU_ADDER_A0 VDD 2.22fF
C476 VDD enable_2/2_input_AND_1/w_n12_9# 0.06fF
C477 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_53_n17# 0.03fF
C478 OUTPUT_ALU_ADDER_B2 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# 0.09fF
C479 ADD_SUB_M OUTPUT_ALU_ADDER_B1 0.47fF
C480 adder_subtractor_0/B0_XOR adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C481 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_A1 0.08fF
C482 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/B0_XOR 0.03fF
C483 comparator_equal_0/A3_B3NOT comparator_equal_0/A3B3 0.15fF
C484 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 1.20fF
C485 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C486 OUTPUT_ALU_ADDER_A3 enable_2/2_input_AND_3/w_35_9# 0.03fF
C487 comparator_equal_0/XNOR_2/OUT comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C488 VDD comparator_equal_0/q1a_NOT_5/w_n12_4# 0.08fF
C489 VDD adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# 0.06fF
C490 and_block_0/2_input_AND_1/w_n12_9# VDD 0.06fF
C491 comparator_equal_0/A3B3 OUTPUT_ALU_COMPARATOR_B1 0.74fF
C492 comparator_equal_0/4_input_AND_2/w_n22_4# comparator_equal_0/4_input_AND_2/OUT 0.09fF
C493 adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/AXORB 0.18fF
C494 adder_subtractor_0/full_adder_0/2_input_AND_0/w_35_9# adder_subtractor_0/full_adder_0/2_input_AND_0/OUT 0.08fF
C495 adder_subtractor_0/B0_XOR OUTPUT_ALU_ADDER_A0 0.75fF
C496 VDD OUTPUT_ALU_ADDER_B1 0.75fF
C497 adder_subtractor_0/full_adder_2/2_input_OR_0/A adder_subtractor_0/full_adder_2/2_input_AND_1/w_35_9# 0.03fF
C498 adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# adder_subtractor_0/B2_XOR 0.07fF
C499 VDD comparator_equal_0/A1B1 1.48fF
C500 GND comparator_equal_0/A3NOT_B3 0.11fF
C501 S0BAR_S1_DECODER enable_1/2_input_AND_0/OUT 0.12fF
C502 adder_subtractor_0/B2_XOR adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# 0.03fF
C503 2_input_AND_0/OUT COMPARATOR_OUT_A_EQUAL_B 0.12fF
C504 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_B0 0.90fF
C505 adder_subtractor_0/B1_XOR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# 0.03fF
C506 GND adder_subtractor_0/full_adder_2/AXORB 0.33fF
C507 GND adder_subtractor_0/full_adder_0/2_input_AND_1/OUT 0.04fF
C508 S0BAR_S1_DECODER OUTPUT_ALU_COMPARATOR_A2 0.25fF
C509 INPUT_ALU_A1 INPUT_ALU_B2 0.59fF
C510 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C511 enable_2/enable enable_2/2_input_AND_6/OUT 0.12fF
C512 OUTPUT_ALU_ADDER_A2 enable_2/2_input_AND_2/OUT 0.05fF
C513 enable_1/2_input_AND_1/w_n12_9# INPUT_ALU_A1 0.07fF
C514 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C515 comparator_equal_0/A1B1 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.58fF
C516 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# comparator_equal_0/A2B2 0.07fF
C517 enable_2/2_input_AND_2/w_n12_9# INPUT_ALU_A2 0.07fF
C518 VDD adder_subtractor_0/full_adder_2/2_input_OR_0/A 0.18fF
C519 adder_subtractor_0/full_adder_0/2_input_OR_0/B VDD 0.12fF
C520 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/4_input_AND_1/w_n22_4# 0.07fF
C521 VDD enable_0/2_input_AND_6/OUT 0.06fF
C522 OUTPUT_ALU_ADDER_B0 OUTPUT_ALU_ADDER_A2 0.25fF
C523 OUTPUT_ALU_ADDER_A0 OUTPUT_ALU_ADDER_B0 0.38fF
C524 VDD adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C525 GND comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C526 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A2B2 0.17fF
C527 OUTPUT_ALU_ADDER_B2 enable_2/2_input_AND_6/w_35_9# 0.12fF
C528 GND OUTPUT_ALU_ADDER_B2 1.53fF
C529 and_block_0/2_input_AND_2/OUT OUTPUT_ALU_ANDBLOCK_B2 0.12fF
C530 OUTPUT_ALU_ANDBLOCK_A1 INPUT_ALU_A2 0.01fF
C531 OUTPUT_ALU_ADDER_A1 INPUT_ALU_A2 0.01fF
C532 enable_1/2_input_AND_4/w_n12_9# enable_1/2_input_AND_4/OUT 0.03fF
C533 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR 0.09fF
C534 VDD enable_1/2_input_AND_1/OUT 0.06fF
C535 GND adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR 0.24fF
C536 VDD adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# 0.03fF
C537 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR 0.09fF
C538 VDD decoder_0/q1a_NOT_1/w_n12_4# 0.05fF
C539 enable_0/2_input_AND_7/w_35_9# enable_0/2_input_AND_7/OUT 0.08fF
C540 and_block_0/2_input_AND_0/w_n12_9# VDD 0.06fF
C541 comparator_equal_0/4_input_AND_1/w_n22_4# comparator_equal_0/A3B3 0.07fF
C542 adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.03fF
C543 adder_subtractor_0/full_adder_1/2_input_OR_0/A adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.05fF
C544 enable_1/2_input_AND_4/w_n12_9# INPUT_ALU_B0 0.07fF
C545 VDD 2_input_OR_0/OUT 0.02fF
C546 OUTPUT_ALU_ADDER_A0 enable_2/2_input_AND_0/OUT 0.05fF
C547 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.08fF
C548 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# comparator_equal_0/A3B3 0.09fF
C549 GND adder_subtractor_0/full_adder_0/2_input_AND_0/OUT 0.04fF
C550 INPUT_ALU_A1 INPUT_ALU_B1 0.55fF
C551 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/A3B3 0.12fF
C552 comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/A2B2 0.09fF
C553 enable_2/enable enable_2/2_input_AND_5/OUT 0.12fF
C554 GND adder_subtractor_0/B2_XOR 0.93fF
C555 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_2/AXORB 0.24fF
C556 comparator_equal_0/q1a_NOT_5/in comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.21fF
C557 enable_2/2_input_AND_1/w_n12_9# enable_2/2_input_AND_1/OUT 0.03fF
C558 VDD comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C559 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A3B3 0.05fF
C560 VDD enable_1/2_input_AND_0/OUT 0.06fF
C561 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_12_2# VDD 0.03fF
C562 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_12_2# 0.03fF
C563 INPUT_ALU_B0 OUTPUT_ALU_COMPARATOR_A3 0.07fF
C564 decoder_0/2_input_AND_3/w_n12_9# S1_DECODER 0.07fF
C565 VDD enable_0/2_input_AND_5/OUT 0.06fF
C566 VDD comparator_equal_0/q1a_NOT_4/w_n12_4# 0.08fF
C567 VDD comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C568 comparator_equal_0/3_input_AND_1/w_n19_2# OUTPUT_ALU_COMPARATOR_B2 0.08fF
C569 VDD comparator_equal_0/3_input_AND_0/OUT 0.09fF
C570 VDD OUTPUT_ALU_COMPARATOR_A2 1.10fF
C571 comparator_equal_0/q1a_NOT_5/w_n12_4# comparator_equal_0/q1a_NOT_5/in 0.12fF
C572 OUTPUT_ALU_ADDER_B1 INPUT_ALU_B2 0.05fF
C573 GND OUTPUT_ALU_COMPARATOR_B0 2.12fF
C574 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_12_2# adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR 0.03fF
C575 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_n34_1# adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.03fF
C576 VDD comparator_equal_0/q1a_NOT_0/w_n12_4# 0.07fF
C577 GND OUTPUT_ALU_COMPARATOR_A0 0.45fF
C578 VDD comparator_equal_0/XNOR_2/w_181_105# 0.06fF
C579 and_block_0/2_input_AND_3/w_n12_9# and_block_0/2_input_AND_3/OUT 0.03fF
C580 adder_subtractor_0/full_adder_0/2_input_OR_0/A adder_subtractor_0/full_adder_0/2_input_OR_0/B 0.45fF
C581 adder_subtractor_0/full_adder_0/2_input_OR_0/w_30_15# adder_subtractor_0/full_adder_0/2_input_OR_0/OUT 0.06fF
C582 VDD decoder_0/2_input_AND_3/w_35_9# 0.03fF
C583 comparator_equal_0/B3_NOT comparator_equal_0/q1a_NOT_0/w_n12_4# 0.04fF
C584 enable_1/2_input_AND_2/w_35_9# enable_1/2_input_AND_2/OUT 0.08fF
C585 adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_AND_0/w_35_9# 0.03fF
C586 adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_2/2_input_OR_0/B 0.07fF
C587 GND OUTPUT_ALU_COMPARATOR_B2 1.61fF
C588 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_S1 0.03fF
C589 VDD adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C590 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C591 enable_0/2_input_AND_6/w_35_9# OUTPUT_ALU_ANDBLOCK_B2 0.07fF
C592 enable_0/2_input_AND_2/w_n12_9# S0_S1_DECODER 0.07fF
C593 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_3/w_n34_1# 0.08fF
C594 GND adder_subtractor_0/full_adder_2/2_input_OR_0/B 0.16fF
C595 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT GND 0.15fF
C596 INPUT_ALU_A1 INPUT_ALU_B0 0.54fF
C597 enable_2/enable enable_2/2_input_AND_4/OUT 0.12fF
C598 enable_1/2_input_AND_3/OUT OUTPUT_ALU_COMPARATOR_A3 0.05fF
C599 comparator_equal_0/A3_B3NOT OUTPUT_ALU_COMPARATOR_B3 0.15fF
C600 GND comparator_equal_0/B1_NOT 0.23fF
C601 enable_2/2_input_AND_6/w_35_9# enable_2/2_input_AND_6/OUT 0.08fF
C602 GND enable_2/2_input_AND_6/OUT 0.04fF
C603 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_53_n17# 0.09fF
C604 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C605 OUTPUT_ALU_COMPARATOR_B1 OUTPUT_ALU_COMPARATOR_B3 0.33fF
C606 VDD enable_0/2_input_AND_4/OUT 0.06fF
C607 enable_1/2_input_AND_1/w_n12_9# enable_1/2_input_AND_1/OUT 0.03fF
C608 S0_S1_DECODER INPUT_ALU_A1 0.68fF
C609 VDD comparator_equal_0/q1a_NOT_3/w_n12_4# 0.07fF
C610 decoder_0/2_input_AND_3/OUT decoder_0/2_input_AND_3/w_n12_9# 0.03fF
C611 enable_1/2_input_AND_3/w_n12_9# enable_1/2_input_AND_3/OUT 0.03fF
C612 VDD adder_subtractor_0/q1d_2_INPUT_XOR_3/w_n34_1# 0.03fF
C613 and_block_0/2_input_AND_1/OUT OUTPUT_ALU_ANDBLOCK_B1 0.12fF
C614 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# comparator_equal_0/B0_NOT 0.07fF
C615 and_block_0/2_input_AND_3/OUT OUTPUT_ALU_ANDBLOCK_B3 0.12fF
C616 comparator_equal_0/A3NOT_B3 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 0.09fF
C617 GND ADDER_SUB_C4 0.16fF
C618 adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_0/AXORB 0.07fF
C619 VDD adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR 0.03fF
C620 comparator_equal_0/B0_NOT comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.08fF
C621 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/full_adder_0/AXORB 0.03fF
C622 comparator_equal_0/B2_NOT OUTPUT_ALU_COMPARATOR_B2 0.04fF
C623 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A3B3 0.15fF
C624 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.09fF
C625 enable_1/2_input_AND_3/w_n12_9# INPUT_ALU_A3 0.07fF
C626 GND enable_1/2_input_AND_7/OUT 0.04fF
C627 adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_3/2_input_OR_0/OUT 0.03fF
C628 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# 0.08fF
C629 VDD enable_0/2_input_AND_3/w_n12_9# 0.06fF
C630 2_input_OR_0/OUT S0BAR_S1BAR_DECODER 0.20fF
C631 S1_DECODER S0_DECODER 0.64fF
C632 INPUT_ALU_A1 INPUT_ALU_A3 0.95fF
C633 enable_2/enable enable_2/2_input_AND_3/OUT 0.12fF
C634 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT ADDER_SUB_C4 0.05fF
C635 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C636 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_12_2# adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C637 OUTPUT_ALU_ANDBLOCK_B2 INPUT_ALU_B3 0.08fF
C638 VDD adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# 0.06fF
C639 adder_subtractor_0/full_adder_0/2_input_AND_1/w_35_9# VDD 0.03fF
C640 VDD enable_2/enable 0.03fF
C641 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# OUTPUT_ALU_COMPARATOR_B1 0.08fF
C642 GND enable_2/2_input_AND_5/OUT 0.04fF
C643 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_12_2# VDD 0.03fF
C644 GND S0_DECODER 0.25fF
C645 VDD enable_0/2_input_AND_3/OUT 0.06fF
C646 OUTPUT_ALU_ANDBLOCK_A1 enable_0/2_input_AND_1/w_35_9# 0.03fF
C647 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C648 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_COMPARATOR_B1 0.08fF
C649 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR VDD 0.03fF
C650 comparator_equal_0/q1a_NOT_5/in OUTPUT_ALU_COMPARATOR_A2 0.72fF
C651 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR 0.09fF
C652 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/full_adder_3/AXORB 0.03fF
C653 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_1/AXORB 0.04fF
C654 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/A3B3 0.29fF
C655 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/4_input_AND_2/w_40_5# 0.03fF
C656 enable_0/2_input_AND_2/w_n12_9# INPUT_ALU_A2 0.07fF
C657 2_input_OR_0/OUT INPUT_ALU_B1 0.18fF
C658 S0BAR_S1_DECODER S1_DECODER 0.17fF
C659 2_input_AND_0/w_n12_9# 2_input_AND_0/OUT 0.03fF
C660 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_n34_1# VDD 0.03fF
C661 adder_subtractor_0/B3_XOR adder_subtractor_0/q1d_2_INPUT_XOR_3/w_53_n17# 0.04fF
C662 GND adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR 0.27fF
C663 adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.03fF
C664 comparator_equal_0/XNOR_0/OUT comparator_equal_0/XNOR_0/w_181_105# 0.13fF
C665 OUTPUT_ALU_ADDER_B2 adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR 0.03fF
C666 adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# ADDER_SUB_C3 0.07fF
C667 and_block_0/2_input_AND_2/w_n12_9# and_block_0/2_input_AND_2/OUT 0.03fF
C668 OUTPUT_ALU_ADDER_A0 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 4.56fF
C669 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_52_34# adder_subtractor_0/full_adder_1/AXORB 0.03fF
C670 S0BAR_S1_DECODER decoder_0/2_input_AND_2/OUT 0.05fF
C671 VDD comparator_equal_0/2_input_AND_0/w_35_9# 0.03fF
C672 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# 0.03fF
C673 VDD adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.06fF
C674 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_ADDER_A0 0.03fF
C675 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_S2 0.03fF
C676 2_input_AND_0/OUT 2_input_AND_0/w_35_9# 0.08fF
C677 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_3/OUT 0.04fF
C678 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C679 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C680 comparator_equal_0/XNOR_0/w_181_105# comparator_equal_0/A0B0 0.06fF
C681 GND S0BAR_S1_DECODER 3.70fF
C682 VDD comparator_equal_0/A2_B2NOT_A3B3XNOR 0.06fF
C683 enable_0/2_input_AND_5/w_35_9# OUTPUT_ALU_ANDBLOCK_B1 0.03fF
C684 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B0_XOR 0.08fF
C685 ADDER_SUB_S0 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR 0.19fF
C686 INPUT_ALU_A1 INPUT_ALU_A2 0.84fF
C687 enable_2/enable enable_2/2_input_AND_2/OUT 0.12fF
C688 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A3B3 0.53fF
C689 OUTPUT_ALU_ADDER_A1 comparator_equal_0/A2NOT_B2_A3B3XNOR 0.19fF
C690 VDD decoder_0/2_input_AND_0/w_35_9# 0.03fF
C691 VDD enable_2/2_input_AND_0/w_35_9# 0.03fF
C692 OUTPUT_ALU_ANDBLOCK_A2 enable_0/2_input_AND_2/OUT 0.05fF
C693 VDD adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# 0.06fF
C694 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_53_n17# 0.03fF
C695 adder_subtractor_0/full_adder_0/2_input_AND_0/w_35_9# VDD 0.03fF
C696 VDD comparator_equal_0/A1NOT 0.10fF
C697 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C698 VDD adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# 0.08fF
C699 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# comparator_equal_0/XNOR_2/OUT 0.03fF
C700 enable_2/2_input_AND_5/w_35_9# enable_2/2_input_AND_5/OUT 0.08fF
C701 GND enable_2/2_input_AND_4/OUT 0.04fF
C702 comparator_equal_0/A0B0 OUTPUT_ALU_COMPARATOR_B1 0.28fF
C703 comparator_equal_0/A3_B3NOT comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.10fF
C704 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 1.54fF
C705 OUTPUT_ALU_ANDBLOCK_A3 OUTPUT_ALU_ANDBLOCK_B2 0.18fF
C706 VDD adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C707 S0_S1_DECODER enable_0/2_input_AND_6/OUT 0.12fF
C708 GND adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.21fF
C709 AND_OUTPUT_A3B3 GND 0.05fF
C710 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR OUTPUT_ALU_COMPARATOR_B1 0.26fF
C711 comparator_equal_0/4_input_AND_2/w_n22_4# OUTPUT_ALU_COMPARATOR_B1 0.08fF
C712 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.17fF
C713 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/B3_XOR 0.03fF
C714 GND comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C715 and_block_0/2_input_AND_0/OUT OUTPUT_ALU_ANDBLOCK_B0 0.12fF
C716 adder_subtractor_0/full_adder_0/2_input_OR_0/A adder_subtractor_0/full_adder_0/2_input_AND_1/w_35_9# 0.03fF
C717 adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# OUTPUT_ALU_ADDER_A0 0.07fF
C718 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR 0.09fF
C719 OUTPUT_ALU_ADDER_B2 OUTPUT_ALU_ADDER_A3 0.33fF
C720 VDD adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.06fF
C721 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_ADDER_A2 0.09fF
C722 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_n34_1# VDD 0.03fF
C723 comparator_equal_0/A1NOT comparator_equal_0/4_input_AND_2/OUT 0.14fF
C724 INPUT_ALU_A1 INPUT_ALU_A0 0.47fF
C725 enable_2/enable enable_2/2_input_AND_0/OUT 0.12fF
C726 enable_1/2_input_AND_0/w_n12_9# enable_1/2_input_AND_0/OUT 0.03fF
C727 GND ADD_SUB_M 1.74fF
C728 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/q1a_NOT_4/out 1.40fF
C729 enable_2/enable INPUT_ALU_B2 0.73fF
C730 adder_subtractor_0/B1_XOR adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR 0.19fF
C731 VDD comparator_equal_0/3_input_AND_1/w_n19_2# 0.06fF
C732 enable_2/enable enable_2/2_input_AND_1/OUT 0.12fF
C733 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C734 VDD adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# 0.03fF
C735 adder_subtractor_0/full_adder_0/2_input_OR_0/w_30_15# VDD 0.03fF
C736 VDD decoder_0/2_input_AND_2/OUT 0.06fF
C737 GND enable_2/2_input_AND_3/OUT 0.04fF
C738 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C739 OUTPUT_ALU_ADDER_A2 adder_subtractor_0/B3_XOR 0.37fF
C740 VDD enable_2/2_input_AND_0/w_n12_9# 0.06fF
C741 adder_subtractor_0/B1_XOR adder_subtractor_0/B2_XOR 0.97fF
C742 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT ADDER_SUB_C2 0.05fF
C743 comparator_equal_0/A1B1 OUTPUT_ALU_COMPARATOR_B1 0.71fF
C744 comparator_equal_0/A0NOT comparator_equal_0/A3B3 0.08fF
C745 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/A2B2 0.08fF
C746 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/A2B2 0.08fF
C747 VDD enable_2/2_input_AND_6/w_35_9# 0.03fF
C748 GND VDD 9.81fF
C749 OUTPUT_ALU_ANDBLOCK_A3 OUTPUT_ALU_ANDBLOCK_B1 0.19fF
C750 OUTPUT_ALU_ANDBLOCK_A2 OUTPUT_ALU_ANDBLOCK_B2 0.52fF
C751 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_12_2# OUTPUT_ALU_ADDER_B1 0.08fF
C752 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_52_34# ADD_SUB_M 0.09fF
C753 VDD comparator_equal_0/q1b_5_INPUT_AND_0/w_50_10# 0.06fF
C754 S0_S1_DECODER enable_0/2_input_AND_5/OUT 0.12fF
C755 GND comparator_equal_0/B3_NOT 0.15fF
C756 enable_2/enable enable_2/2_input_AND_7/OUT 0.12fF
C757 AND_OUTPUT_A2B2 GND 0.05fF
C758 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/A2B2 2.19fF
C759 comparator_equal_0/A2NOT comparator_equal_0/A3B3 0.01fF
C760 enable_0/2_input_AND_7/w_n12_9# enable_0/2_input_AND_7/OUT 0.03fF
C761 adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.03fF
C762 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/4_input_AND_1/w_40_5# 0.03fF
C763 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/q1a_NOT_4/out 0.04fF
C764 adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# OUTPUT_ALU_ADDER_A3 0.07fF
C765 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_52_34# adder_subtractor_0/full_adder_2/AXORB 0.03fF
C766 and_block_0/2_input_AND_1/w_n12_9# and_block_0/2_input_AND_1/OUT 0.03fF
C767 GND comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.06fF
C768 decoder_0/2_input_AND_0/w_35_9# decoder_0/2_input_AND_0/OUT 0.08fF
C769 OUTPUT_ALU_ANDBLOCK_A0 enable_0/2_input_AND_0/OUT 0.05fF
C770 VDD adder_subtractor_0/full_adder_3/2_input_OR_0/OUT 0.02fF
C771 enable_2/2_input_AND_0/w_35_9# enable_2/2_input_AND_0/OUT 0.08fF
C772 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# OUTPUT_ALU_COMPARATOR_B0 0.07fF
C773 enable_1/2_input_AND_0/w_35_9# enable_1/2_input_AND_0/OUT 0.08fF
C774 comparator_equal_0/B1_NOT comparator_equal_0/A2B2 1.02fF
C775 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR ADDER_SUB_C2 0.03fF
C776 ADDER_SUB_S2 adder_subtractor_0/full_adder_2/AXORB 0.18fF
C777 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_0/AXORB 0.24fF
C778 GND adder_subtractor_0/B0_XOR 0.52fF
C779 INPUT_ALU_B3 INPUT_ALU_A1 0.54fF
C780 S0_S1_DECODER decoder_0/2_input_AND_3/w_35_9# 0.03fF
C781 GND comparator_equal_0/4_input_AND_2/OUT 0.11fF
C782 enable_2/enable INPUT_ALU_B1 1.13fF
C783 OUTPUT_ALU_ANDBLOCK_A2 enable_0/2_input_AND_2/w_35_9# 0.03fF
C784 GND COMPARATOR_OUT_A_GREATERTHAN_B 0.05fF
C785 enable_0/2_input_AND_4/w_35_9# OUTPUT_ALU_ANDBLOCK_B0 0.03fF
C786 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.08fF
C787 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.05fF
C788 comparator_equal_0/B0_NOT comparator_equal_0/A3B3 0.08fF
C789 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_12_2# 0.03fF
C790 VDD decoder_0/2_input_AND_3/OUT 0.06fF
C791 decoder_0/2_input_AND_0/w_35_9# S0BAR_S1BAR_DECODER 0.03fF
C792 INPUT_ALU_A3 OUTPUT_ALU_COMPARATOR_A2 0.02fF
C793 enable_2/2_input_AND_4/w_35_9# enable_2/2_input_AND_4/OUT 0.08fF
C794 GND enable_2/2_input_AND_2/OUT 0.04fF
C795 VDD comparator_equal_0/XNOR_3/OUT 0.12fF
C796 VDD comparator_equal_0/B2_NOT 0.10fF
C797 VDD comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C798 VDD enable_2/2_input_AND_5/w_35_9# 0.03fF
C799 OUTPUT_ALU_ANDBLOCK_A3 OUTPUT_ALU_ANDBLOCK_B0 0.19fF
C800 OUTPUT_ALU_ANDBLOCK_A2 OUTPUT_ALU_ANDBLOCK_B1 0.17fF
C801 enable_0/2_input_AND_2/OUT enable_0/2_input_AND_2/w_35_9# 0.08fF
C802 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C803 enable_1/2_input_AND_6/w_35_9# OUTPUT_ALU_COMPARATOR_B2 0.12fF
C804 S0_S1_DECODER enable_0/2_input_AND_4/OUT 0.12fF
C805 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_12_2# OUTPUT_ALU_ADDER_B3 0.08fF
C806 GND OUTPUT_ALU_ADDER_B0 1.09fF
C807 GND enable_0/2_input_AND_1/OUT 0.04fF
C808 AND_OUTPUT_A1B1 GND 0.05fF
C809 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/3_input_AND_1/OUT 0.08fF
C810 VDD comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C811 and_block_0/2_input_AND_3/w_n12_9# OUTPUT_ALU_ANDBLOCK_A3 0.07fF
C812 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# comparator_equal_0/A1B1 0.07fF
C813 OUTPUT_ALU_COMPARATOR_A1 OUTPUT_ALU_COMPARATOR_B3 0.27fF
C814 comparator_equal_0/3_input_AND_0/w_n19_2# comparator_equal_0/A3B3 0.08fF
C815 adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_AND_0/w_35_9# 0.03fF
C816 adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_0/2_input_OR_0/B 0.07fF
C817 OUTPUT_ALU_ADDER_B3 adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.08fF
C818 VDD comparator_equal_0/2_input_AND_1/w_n12_9# 0.06fF
C819 GND enable_1/2_input_AND_6/OUT 0.04fF
C820 enable_0/2_input_AND_6/w_35_9# enable_0/2_input_AND_6/OUT 0.08fF
C821 comparator_equal_0/A3B3 comparator_equal_0/XNOR_3/w_181_105# 0.06fF
C822 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A1B1 0.08fF
C823 adder_subtractor_0/full_adder_0/2_input_OR_0/A GND 0.44fF
C824 enable_2/enable INPUT_ALU_B0 0.64fF
C825 enable_1/2_input_AND_2/OUT OUTPUT_ALU_COMPARATOR_A2 0.05fF
C826 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR ADDER_SUB_C3 0.51fF
C827 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_2/AXORB 0.19fF
C828 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR 0.09fF
C829 enable_2/2_input_AND_0/w_n12_9# enable_2/2_input_AND_0/OUT 0.03fF
C830 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_12_2# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C831 GND decoder_0/2_input_AND_0/OUT 0.04fF
C832 S0_S1_DECODER enable_0/2_input_AND_3/w_n12_9# 0.07fF
C833 GND enable_2/2_input_AND_0/OUT 0.04fF
C834 VDD enable_2/2_input_AND_7/w_n12_9# 0.07fF
C835 VDD comparator_equal_0/4_input_AND_0/w_n22_4# 0.05fF
C836 GND INPUT_ALU_B2 1.94fF
C837 ADD_SUB_M OUTPUT_ALU_ADDER_B3 0.88fF
C838 comparator_equal_0/A3B3 OUTPUT_ALU_COMPARATOR_B3 0.53fF
C839 GND enable_2/2_input_AND_1/OUT 0.04fF
C840 comparator_equal_0/B1_NOT comparator_equal_0/4_input_AND_1/OUT 0.09fF
C841 VDD enable_0/2_input_AND_7/OUT 0.06fF
C842 GND comparator_equal_0/q1a_NOT_5/in 0.04fF
C843 VDD enable_2/2_input_AND_4/w_35_9# 0.03fF
C844 OUTPUT_ALU_ANDBLOCK_A2 OUTPUT_ALU_ANDBLOCK_B0 0.17fF
C845 OUTPUT_ALU_ANDBLOCK_A3 OUTPUT_ALU_ANDBLOCK_B3 0.55fF
C846 OUTPUT_ALU_ANDBLOCK_A1 OUTPUT_ALU_ANDBLOCK_B1 0.50fF
C847 OUTPUT_ALU_COMPARATOR_A1 OUTPUT_ALU_COMPARATOR_A3 0.22fF
C848 GND S0BAR_S1BAR_DECODER 0.05fF
C849 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 0.10fF
C850 GND decoder_0/2_input_AND_1/OUT 0.04fF
C851 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A0B0 0.14fF
C852 S0_S1_DECODER enable_0/2_input_AND_3/OUT 0.12fF
C853 VDD OUTPUT_ALU_ADDER_B3 0.50fF
C854 enable_0/2_input_AND_3/w_n12_9# INPUT_ALU_A3 0.07fF
C855 AND_OUTPUT_A0B0 GND 0.05fF
C856 OUTPUT_ALU_ANDBLOCK_A3 enable_0/2_input_AND_3/w_35_9# 0.12fF
C857 adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_1/2_input_OR_0/OUT 0.03fF
C858 comparator_equal_0/q1c_4_INPUT_OR_1/w_41_n9# comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.10fF
C859 enable_1/2_input_AND_2/w_n12_9# S0BAR_S1_DECODER 0.07fF
C860 adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_3/2_input_OR_0/A 0.07fF
C861 decoder_0/A0_BAR S1_DECODER 0.59fF
C862 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# 0.09fF
C863 GND enable_2/2_input_AND_7/OUT 0.04fF
C864 VDD enable_0/2_input_AND_1/w_n12_9# 0.06fF
C865 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/2_input_AND_0/w_n12_9# 0.07fF
C866 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_n34_1# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C867 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C868 GND enable_1/2_input_AND_5/OUT 0.04fF
C869 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B2_XOR 0.11fF
C870 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A3B3 0.29fF
C871 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/OUT 0.15fF
C872 VDD comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C873 enable_2/enable INPUT_ALU_A3 0.61fF
C874 and_block_0/2_input_AND_0/w_n12_9# and_block_0/2_input_AND_0/OUT 0.03fF
C875 VDD enable_2/2_input_AND_7/w_35_9# 0.03fF
C876 GND decoder_0/A0_BAR 0.41fF
C877 GND comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C878 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# OUTPUT_ALU_COMPARATOR_B1 0.09fF
C879 GND INPUT_ALU_B1 2.36fF
C880 decoder_0/A1_BAR decoder_0/2_input_AND_1/w_n12_9# 0.07fF
C881 enable_1/2_input_AND_4/w_35_9# OUTPUT_ALU_COMPARATOR_B0 0.12fF
C882 enable_0/2_input_AND_2/OUT enable_0/2_input_AND_2/w_n12_9# 0.03fF
C883 enable_2/2_input_AND_3/w_35_9# enable_2/2_input_AND_3/OUT 0.08fF
C884 enable_1/2_input_AND_7/w_n12_9# enable_1/2_input_AND_7/OUT 0.03fF
C885 comparator_equal_0/XNOR_1/OUT OUTPUT_ALU_COMPARATOR_B1 0.15fF
C886 VDD enable_2/2_input_AND_3/w_35_9# 0.03fF
C887 OUTPUT_ALU_ANDBLOCK_A1 OUTPUT_ALU_ANDBLOCK_B0 0.19fF
C888 INPUT_ALU_A0 decoder_0/2_input_AND_3/w_35_9# 0.02fF
C889 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# 0.03fF
C890 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/full_adder_1/AXORB 0.03fF
C891 comparator_equal_0/A1B1 comparator_equal_0/4_input_AND_0/OUT 0.09fF
C892 enable_1/2_input_AND_7/OUT enable_1/2_input_AND_7/w_35_9# 0.08fF
C893 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_3/AXORB 0.19fF
C894 OUTPUT_ALU_ADDER_B0 enable_2/2_input_AND_4/w_35_9# 0.03fF
C895 GND ADDER_SUB_S3 0.05fF
C896 GND adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR 0.04fF
C897 GND comparator_equal_0/2_input_AND_1/OUT 0.04fF
C898 comparator_equal_0/XNOR_0/OUT comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C899 VDD adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR 0.03fF
C900 adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# ADDER_SUB_C1 0.07fF
C901 and_block_0/2_input_AND_2/w_n12_9# OUTPUT_ALU_ANDBLOCK_A2 0.07fF
C902 OUTPUT_ALU_ADDER_A0 comparator_equal_0/A2NOT_B2_A3B3XNOR 0.30fF
C903 VDD ADDER_SUB_C3 0.15fF
C904 VDD adder_subtractor_0/full_adder_1/AXORB 0.43fF
C905 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/4_input_AND_2/OUT 0.04fF
C906 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A0B0 0.38fF
C907 GND enable_1/2_input_AND_4/OUT 0.04fF
C908 adder_subtractor_0/full_adder_3/AXORB adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.12fF
C909 adder_subtractor_0/B2_XOR adder_subtractor_0/full_adder_2/AXORB 0.18fF
C910 VDD comparator_equal_0/q1c_4_INPUT_OR_0/w_41_n9# 0.09fF
C911 enable_0/2_input_AND_5/w_35_9# enable_0/2_input_AND_5/OUT 0.08fF
C912 VDD comparator_equal_0/2_input_AND_0/OUT 0.06fF
C913 enable_0/2_input_AND_1/OUT enable_0/2_input_AND_1/w_n12_9# 0.03fF
C914 VDD adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# 0.10fF
C915 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_12_2# OUTPUT_ALU_ADDER_A2 0.08fF
C916 enable_2/enable INPUT_ALU_A2 0.76fF
C917 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C918 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.19fF
C919 ADDER_SUB_C4 adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.08fF
C920 comparator_equal_0/A3_B3NOT comparator_equal_0/2_input_AND_0/w_35_9# 0.03fF
C921 adder_subtractor_0/B2_XOR adder_subtractor_0/q1d_2_INPUT_XOR_2/w_53_n17# 0.04fF
C922 VDD comparator_equal_0/A2B2 1.39fF
C923 comparator_equal_0/A1B1 comparator_equal_0/XNOR_1/w_181_105# 0.06fF
C924 GND COMPARATOR_OUT_A_EQUAL_B 0.11fF
C925 VDD enable_1/2_input_AND_2/w_n12_9# 0.06fF
C926 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# OUTPUT_ALU_COMPARATOR_A2 0.08fF
C927 GND INPUT_ALU_B0 2.48fF
C928 ADD_SUB_M OUTPUT_ALU_ADDER_A3 0.46fF
C929 ADD_SUB_M adder_subtractor_0/B1_XOR 0.18fF
C930 VDD adder_subtractor_0/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C931 comparator_equal_0/A3_B3NOT comparator_equal_0/A2_B2NOT_A3B3XNOR 2.07fF
C932 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.10fF
C933 comparator_equal_0/A0B0 comparator_equal_0/A3B3 0.34fF
C934 adder_subtractor_0/B2_XOR OUTPUT_ALU_ADDER_B2 0.27fF
C935 comparator_equal_0/3_input_AND_0/a_n3_n34# OUTPUT_ALU_COMPARATOR_A2 0.01fF
C936 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C937 VDD enable_2/2_input_AND_2/w_35_9# 0.03fF
C938 decoder_0/A1_BAR S0_DECODER 0.57fF
C939 S0BAR_S1_DECODER enable_1/2_input_AND_7/w_n12_9# 0.07fF
C940 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/B1_XOR 0.03fF
C941 comparator_equal_0/4_input_AND_2/w_n22_4# comparator_equal_0/A3B3 0.28fF
C942 enable_2/2_input_AND_7/w_n12_9# enable_2/2_input_AND_7/OUT 0.03fF
C943 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B3_XOR 0.11fF
C944 and_block_0/2_input_AND_3/OUT GND 0.04fF
C945 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/A2B2 0.74fF
C946 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/A3B3 0.22fF
C947 comparator_equal_0/q1c_4_INPUT_OR_0/w_41_n9# COMPARATOR_OUT_A_GREATERTHAN_B 0.05fF
C948 comparator_equal_0/A3_B3NOT comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.09fF
C949 comparator_equal_0/q1a_NOT_4/w_n12_4# comparator_equal_0/q1a_NOT_4/out 0.04fF
C950 GND S0_S1_DECODER 3.35fF
C951 OUTPUT_ALU_ANDBLOCK_A0 OUTPUT_ALU_ANDBLOCK_B0 0.44fF
C952 OUTPUT_ALU_ADDER_A3 enable_2/2_input_AND_3/OUT 0.05fF
C953 VDD comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# 0.15fF
C954 VDD OUTPUT_ALU_ADDER_A3 1.05fF
C955 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_n34_1# adder_subtractor_0/B2_XOR 0.08fF
C956 VDD adder_subtractor_0/B1_XOR 0.67fF
C957 comparator_equal_0/A2B2 comparator_equal_0/4_input_AND_2/OUT 0.09fF
C958 OUTPUT_ALU_COMPARATOR_B1 comparator_equal_0/A1NOT 0.67fF
C959 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A1B1 0.36fF
C960 enable_2/enable INPUT_ALU_A0 0.74fF
C961 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C962 GND enable_1/2_input_AND_3/OUT 0.04fF
C963 adder_subtractor_0/full_adder_2/2_input_OR_0/A adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.05fF
C964 enable_2/enable enable_2/2_input_AND_6/w_n12_9# 0.07fF
C965 ADDER_SUB_CFINAL adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.19fF
C966 S0BAR_S1_DECODER decoder_0/2_input_AND_2/w_35_9# 0.03fF
C967 GND comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.14fF
C968 VDD comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.32fF
C969 VDD enable_1/2_input_AND_6/w_35_9# 0.03fF
C970 OUTPUT_ALU_ADDER_B3 enable_2/2_input_AND_7/OUT 0.05fF
C971 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_12_2# 0.03fF
C972 GND adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C973 comparator_equal_0/2_input_AND_1/w_n12_9# comparator_equal_0/2_input_AND_1/OUT 0.03fF
C974 VDD comparator_equal_0/3_input_AND_1/OUT 0.09fF
C975 VDD enable_0/2_input_AND_6/w_n12_9# 0.07fF
C976 GND INPUT_ALU_A3 2.14fF
C977 VDD decoder_0/2_input_AND_2/w_n12_9# 0.06fF
C978 comparator_equal_0/A1B1 comparator_equal_0/A3B3 1.84fF
C979 adder_subtractor_0/full_adder_2/2_input_OR_0/w_30_15# ADDER_SUB_C3 0.03fF
C980 enable_2/2_input_AND_2/w_35_9# enable_2/2_input_AND_2/OUT 0.08fF
C981 and_block_0/2_input_AND_2/w_n12_9# OUTPUT_ALU_ANDBLOCK_B2 0.07fF
C982 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_12_2# OUTPUT_ALU_ADDER_B0 0.08fF
C983 OUTPUT_ALU_ANDBLOCK_A0 INPUT_ALU_A1 0.07fF
C984 S0_S1_DECODER decoder_0/2_input_AND_3/OUT 0.05fF
C985 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C986 GND adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.21fF
C987 GND adder_subtractor_0/full_adder_3/AXORB 0.33fF
C988 GND adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.04fF
C989 and_block_0/2_input_AND_2/OUT GND 0.04fF
C990 enable_2/2_input_AND_7/w_35_9# enable_2/2_input_AND_7/OUT 0.08fF
C991 enable_1/2_input_AND_1/OUT OUTPUT_ALU_COMPARATOR_A1 0.05fF
C992 OUTPUT_ALU_ADDER_B2 enable_2/2_input_AND_6/OUT 0.05fF
C993 OUTPUT_ALU_COMPARATOR_A3 OUTPUT_ALU_COMPARATOR_B3 1.29fF
C994 adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# OUTPUT_ALU_ADDER_A1 0.07fF
C995 and_block_0/2_input_AND_1/w_n12_9# OUTPUT_ALU_ANDBLOCK_A1 0.07fF
C996 GND comparator_equal_0/A3_B3NOT 0.11fF
C997 VDD adder_subtractor_0/full_adder_3/2_input_OR_0/A 0.18fF
C998 VDD adder_subtractor_0/full_adder_1/2_input_OR_0/B 0.12fF
C999 OUTPUT_ALU_ADDER_B0 OUTPUT_ALU_ADDER_A3 0.24fF
C1000 OUTPUT_ALU_ADDER_A1 OUTPUT_ALU_ADDER_B1 0.25fF
C1001 INPUT_ALU_A2 S1_DECODER 0.27fF
C1002 VDD enable_1/2_input_AND_7/w_n12_9# 0.07fF
C1003 VDD adder_subtractor_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C1004 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR ADD_SUB_M 0.03fF
C1005 ADDER_SUB_S0 adder_subtractor_0/full_adder_0/AXORB 0.18fF
C1006 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR comparator_equal_0/4_input_AND_1/OUT 0.04fF
C1007 enable_2/enable enable_2/2_input_AND_5/w_n12_9# 0.07fF
C1008 INPUT_ALU_B3 enable_2/enable 0.94fF
C1009 GND enable_1/2_input_AND_2/OUT 0.04fF
C1010 adder_subtractor_0/B3_XOR adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.12fF
C1011 GND OUTPUT_ALU_COMPARATOR_B1 1.85fF
C1012 enable_0/2_input_AND_4/w_35_9# enable_0/2_input_AND_4/OUT 0.08fF
C1013 VDD COMPARATOR_A_EQUAL_B_FINAL 0.02fF
C1014 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_12_2# adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1015 comparator_equal_0/q1a_NOT_5/w_n12_4# comparator_equal_0/A2NOT 0.04fF
C1016 VDD enable_1/2_input_AND_5/w_35_9# 0.03fF
C1017 comparator_equal_0/A1B1 comparator_equal_0/A0NOT 0.08fF
C1018 decoder_0/A1_BAR decoder_0/2_input_AND_0/w_n12_9# 0.07fF
C1019 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_B0 0.64fF
C1020 VDD enable_1/2_input_AND_7/w_35_9# 0.03fF
C1021 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/w_12_2# 0.08fF
C1022 GND adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C1023 comparator_equal_0/q1a_NOT_5/in comparator_equal_0/A2B2 0.31fF
C1024 comparator_equal_0/A3NOT_B3 comparator_equal_0/2_input_AND_1/w_35_9# 0.03fF
C1025 VDD enable_0/2_input_AND_5/w_n12_9# 0.06fF
C1026 GND INPUT_ALU_A2 3.09fF
C1027 VDD comparator_equal_0/3_input_AND_0/w_34_3# 0.03fF
C1028 OUTPUT_ALU_COMPARATOR_B0 OUTPUT_ALU_COMPARATOR_B2 0.06fF
C1029 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_B2 0.84fF
C1030 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.08fF
C1031 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR VDD 0.03fF
C1032 VDD decoder_0/2_input_AND_2/w_35_9# 0.03fF
C1033 OUTPUT_ALU_COMPARATOR_A1 OUTPUT_ALU_COMPARATOR_A2 0.23fF
C1034 VDD decoder_0/A1_BAR 1.20fF
C1035 VDD comparator_equal_0/q1a_NOT_7/w_n12_4# 0.07fF
C1036 enable_1/2_input_AND_6/w_35_9# enable_1/2_input_AND_6/OUT 0.08fF
C1037 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# OUTPUT_ALU_ADDER_B3 0.09fF
C1038 GND adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.04fF
C1039 comparator_equal_0/3_input_AND_1/w_34_3# comparator_equal_0/3_input_AND_1/OUT 0.06fF
C1040 enable_0/2_input_AND_7/OUT S0_S1_DECODER 0.12fF
C1041 GND adder_subtractor_0/B3_XOR 0.79fF
C1042 and_block_0/2_input_AND_1/OUT GND 0.04fF
C1043 VDD comparator_equal_0/XNOR_2/OUT 0.13fF
C1044 VDD adder_subtractor_0/q1d_2_INPUT_XOR_4/w_12_2# 0.03fF
C1045 and_block_0/2_input_AND_3/w_35_9# AND_OUTPUT_A3B3 0.03fF
C1046 VDD adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.03fF
C1047 comparator_equal_0/B0_NOT comparator_equal_0/A1B1 0.73fF
C1048 enable_2/enable enable_2/2_input_AND_4/w_n12_9# 0.07fF
C1049 ADDER_SUB_S3 ADDER_SUB_C3 0.15fF
C1050 adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.05fF
C1051 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR ADDER_SUB_C1 0.51fF
C1052 comparator_equal_0/A0B0 OUTPUT_ALU_COMPARATOR_B3 0.36fF
C1053 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C1054 INPUT_ALU_A0 enable_2/2_input_AND_0/w_n12_9# 0.07fF
C1055 enable_0/2_input_AND_6/w_n12_9# INPUT_ALU_B2 0.07fF
C1056 enable_0/2_input_AND_1/w_n12_9# S0_S1_DECODER 0.07fF
C1057 VDD enable_1/2_input_AND_4/w_35_9# 0.03fF
C1058 GND INPUT_ALU_A0 1.50fF
C1059 VDD enable_0/2_input_AND_7/w_35_9# 0.03fF
C1060 enable_0/2_input_AND_6/OUT OUTPUT_ALU_ANDBLOCK_B2 0.05fF
C1061 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C1062 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR OUTPUT_ALU_COMPARATOR_B3 1.13fF
C1063 comparator_equal_0/XNOR_1/OUT comparator_equal_0/XNOR_1/w_181_105# 0.13fF
C1064 VDD enable_0/2_input_AND_4/w_n12_9# 0.06fF
C1065 comparator_equal_0/4_input_AND_1/w_40_5# comparator_equal_0/q1a_NOT_2/vdd 0.03fF
C1066 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C1067 OUTPUT_ALU_ANDBLOCK_A3 enable_0/2_input_AND_3/OUT 0.05fF
C1068 and_block_0/2_input_AND_1/w_n12_9# OUTPUT_ALU_ANDBLOCK_B1 0.07fF
C1069 and_block_0/2_input_AND_3/w_n12_9# OUTPUT_ALU_ANDBLOCK_B3 0.07fF
C1070 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# comparator_equal_0/A3NOT_B3 0.13fF
C1071 GND comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.06fF
C1072 GND adder_subtractor_0/full_adder_3/2_input_OR_0/B 0.16fF
C1073 GND adder_subtractor_0/full_adder_1/2_input_OR_0/OUT 0.15fF
C1074 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1075 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C1076 comparator_equal_0/q1b_5_INPUT_AND_0/w_50_10# comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.07fF
C1077 and_block_0/2_input_AND_3/w_35_9# VDD 0.03fF
C1078 and_block_0/2_input_AND_0/OUT GND 0.04fF
C1079 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 1.40fF
C1080 adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_1/2_input_OR_0/A 0.07fF
C1081 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A0B0 0.17fF
C1082 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/XNOR_1/OUT 0.18fF
C1083 adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.03fF
C1084 INPUT_ALU_A0 decoder_0/2_input_AND_3/OUT 0.09fF
C1085 decoder_0/2_input_AND_3/w_n12_9# S0_DECODER 0.07fF
C1086 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/q1a_NOT_6/w_n12_4# 0.09fF
C1087 2_input_OR_0/w_n23_15# 2_input_OR_0/OUT 0.03fF
C1088 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_0/AXORB 0.04fF
C1089 enable_2/enable enable_2/2_input_AND_3/w_n12_9# 0.07fF
C1090 adder_subtractor_0/full_adder_3/2_input_OR_0/B adder_subtractor_0/full_adder_3/2_input_OR_0/OUT 0.20fF
C1091 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A2 0.03fF
C1092 and_block_0/2_input_AND_0/w_n12_9# OUTPUT_ALU_ANDBLOCK_A0 0.07fF
C1093 decoder_0/A0_BAR decoder_0/2_input_AND_2/w_n12_9# 0.07fF
C1094 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.47fF
C1095 comparator_equal_0/A1B1 OUTPUT_ALU_COMPARATOR_B3 0.76fF
C1096 VDD enable_1/2_input_AND_3/w_35_9# 0.03fF
C1097 VDD comparator_equal_0/A3NOT_B3 0.02fF
C1098 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C1099 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# comparator_equal_0/XNOR_0/OUT 0.03fF
C1100 2_input_OR_0/OUT 2_input_OR_0/w_30_15# 0.06fF
C1101 GND INPUT_ALU_B3 1.94fF
C1102 GND adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR 0.04fF
C1103 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR GND 0.27fF
C1104 ADD_SUB_M OUTPUT_ALU_ADDER_B2 0.62fF
C1105 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_53_n17# 0.03fF
C1106 VDD adder_subtractor_0/full_adder_2/AXORB 0.43fF
C1107 adder_subtractor_0/full_adder_0/2_input_AND_1/OUT VDD 0.06fF
C1108 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C1109 decoder_0/2_input_AND_1/w_n12_9# S0_DECODER 0.07fF
C1110 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_53_n17# 0.09fF
C1111 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_n34_1# VDD 0.03fF
C1112 GND comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C1113 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_1/AXORB 0.19fF
C1114 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR 0.08fF
C1115 enable_1/2_input_AND_5/w_35_9# enable_1/2_input_AND_5/OUT 0.08fF
C1116 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_53_n17# 0.09fF
C1117 OUTPUT_ALU_ADDER_A3 INPUT_ALU_B0 0.14fF
C1118 GND comparator_equal_0/q1a_NOT_4/out 0.50fF
C1119 decoder_0/A1_BAR S0BAR_S1BAR_DECODER 0.07fF
C1120 VDD comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1121 VDD adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# 0.06fF
C1122 VDD adder_subtractor_0/full_adder_1/2_input_AND_1/w_35_9# 0.03fF
C1123 and_block_0/2_input_AND_2/w_35_9# VDD 0.03fF
C1124 VDD OUTPUT_ALU_ADDER_B2 0.94fF
C1125 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A1B1 0.17fF
C1126 adder_subtractor_0/B3_XOR OUTPUT_ALU_ADDER_B3 0.33fF
C1127 ADDER_SUB_C4 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_52_34# 0.03fF
C1128 OUTPUT_ALU_ADDER_A0 INPUT_ALU_A1 0.04fF
C1129 ADD_SUB_M adder_subtractor_0/B2_XOR 0.18fF
C1130 adder_subtractor_0/full_adder_3/2_input_AND_1/w_35_9# adder_subtractor_0/full_adder_3/2_input_AND_1/OUT 0.08fF
C1131 ADDER_SUB_C3 adder_subtractor_0/full_adder_3/AXORB 0.93fF
C1132 adder_subtractor_0/full_adder_1/AXORB adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.12fF
C1133 OUTPUT_ALU_ADDER_A0 adder_subtractor_0/full_adder_0/AXORB 0.18fF
C1134 and_block_0/2_input_AND_2/w_35_9# AND_OUTPUT_A2B2 0.04fF
C1135 enable_2/2_input_AND_1/w_n12_9# INPUT_ALU_A1 0.07fF
C1136 VDD adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1137 enable_2/enable enable_2/2_input_AND_2/w_n12_9# 0.07fF
C1138 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_53_n17# ADDER_SUB_S2 0.04fF
C1139 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_12_2# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C1140 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1141 enable_0/2_input_AND_5/w_n12_9# INPUT_ALU_B1 0.07fF
C1142 ADDER_SUB_C4 ADDER_SUB_CFINAL 0.18fF
C1143 comparator_equal_0/3_input_AND_0/w_n19_2# comparator_equal_0/3_input_AND_0/OUT 0.06fF
C1144 VDD comparator_equal_0/4_input_AND_2/w_40_5# 0.03fF
C1145 comparator_equal_0/3_input_AND_0/w_n19_2# OUTPUT_ALU_COMPARATOR_A2 0.08fF
C1146 GND comparator_equal_0/4_input_AND_0/OUT 0.11fF
C1147 enable_0/2_input_AND_5/OUT OUTPUT_ALU_ANDBLOCK_B1 0.05fF
C1148 VDD adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C1149 enable_1/2_input_AND_2/w_35_9# OUTPUT_ALU_COMPARATOR_A2 0.13fF
C1150 GND adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C1151 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A1NOT 0.04fF
C1152 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# comparator_equal_0/A2_B2NOT_A3B3XNOR 0.10fF
C1153 decoder_0/A0_BAR decoder_0/A1_BAR 0.55fF
C1154 comparator_equal_0/B2_NOT comparator_equal_0/q1a_NOT_1/w_n12_4# 0.04fF
C1155 comparator_equal_0/A3_B3NOT comparator_equal_0/2_input_AND_0/OUT 0.05fF
C1156 VDD adder_subtractor_0/B2_XOR 1.11fF
C1157 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT VDD 0.06fF
C1158 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# 0.08fF
C1159 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_12_2# OUTPUT_ALU_ADDER_A1 0.08fF
C1160 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_2/OUT 0.04fF
C1161 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1162 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C1163 S0_S1_DECODER enable_0/2_input_AND_6/w_n12_9# 0.07fF
C1164 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/B1_XOR 0.11fF
C1165 OUTPUT_ALU_ANDBLOCK_A3 GND 0.34fF
C1166 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/A3B3 0.75fF
C1167 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.06fF
C1168 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.05fF
C1169 comparator_equal_0/q1a_NOT_3/w_n12_4# comparator_equal_0/B0_NOT 0.04fF
C1170 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C1171 and_block_0/2_input_AND_0/w_n12_9# OUTPUT_ALU_ANDBLOCK_B0 0.07fF
C1172 S0BAR_S1_DECODER enable_1/2_input_AND_7/OUT 0.12fF
C1173 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_52_34# ADDER_SUB_CFINAL 0.03fF
C1174 comparator_equal_0/A3B3 comparator_equal_0/A1NOT 0.05fF
C1175 comparator_equal_0/A2B2 OUTPUT_ALU_COMPARATOR_B1 2.63fF
C1176 comparator_equal_0/4_input_AND_2/w_40_5# comparator_equal_0/4_input_AND_2/OUT 0.07fF
C1177 VDD adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# 0.06fF
C1178 VDD adder_subtractor_0/full_adder_1/2_input_AND_0/w_35_9# 0.03fF
C1179 and_block_0/2_input_AND_1/w_35_9# VDD 0.03fF
C1180 enable_1/2_input_AND_2/w_n12_9# enable_1/2_input_AND_2/OUT 0.03fF
C1181 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/q1a_NOT_0/w_n12_4# 0.10fF
C1182 adder_subtractor_0/full_adder_0/2_input_OR_0/A adder_subtractor_0/full_adder_0/2_input_AND_1/OUT 0.05fF
C1183 INPUT_ALU_B3 enable_2/2_input_AND_7/w_n12_9# 0.07fF
C1184 OUTPUT_ALU_ADDER_A3 adder_subtractor_0/full_adder_3/AXORB 0.15fF
C1185 adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.03fF
C1186 GND comparator_equal_0/A2NOT_B2_A3B3XNOR 0.10fF
C1187 VDD OUTPUT_ALU_COMPARATOR_B0 0.90fF
C1188 VDD decoder_0/2_input_AND_3/w_n12_9# 0.06fF
C1189 VDD OUTPUT_ALU_COMPARATOR_A0 0.68fF
C1190 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR adder_subtractor_0/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C1191 enable_1/2_input_AND_2/w_n12_9# INPUT_ALU_A2 0.07fF
C1192 comparator_equal_0/q1a_NOT_4/out comparator_equal_0/2_input_AND_1/w_n12_9# 0.07fF
C1193 comparator_equal_0/A1B1 comparator_equal_0/A0B0 1.20fF
C1194 GND adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.04fF
C1195 VDD OUTPUT_ALU_COMPARATOR_B2 1.50fF
C1196 GND comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.63fF
C1197 S0BAR_S1_DECODER S0_DECODER 0.02fF
C1198 adder_subtractor_0/full_adder_0/2_input_OR_0/w_30_15# ADDER_SUB_C1 0.03fF
C1199 comparator_equal_0/A1B1 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.33fF
C1200 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/q1a_NOT_4/w_n12_4# 0.09fF
C1201 VDD adder_subtractor_0/full_adder_2/2_input_OR_0/B 0.12fF
C1202 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT VDD 0.02fF
C1203 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C1204 OUTPUT_ALU_COMPARATOR_A3 OUTPUT_ALU_COMPARATOR_A2 0.22fF
C1205 OUTPUT_ALU_ADDER_A2 OUTPUT_ALU_ADDER_B1 0.35fF
C1206 VDD decoder_0/2_input_AND_1/w_n12_9# 0.06fF
C1207 GND OUTPUT_ALU_COMPARATOR_A1 1.54fF
C1208 S0_S1_DECODER enable_0/2_input_AND_5/w_n12_9# 0.07fF
C1209 GND enable_0/2_input_AND_0/OUT 0.04fF
C1210 GND ADDER_SUB_C1 0.81fF
C1211 OUTPUT_ALU_ANDBLOCK_A2 GND 0.32fF
C1212 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR OUTPUT_ALU_COMPARATOR_B2 0.68fF
C1213 comparator_equal_0/3_input_AND_1/w_n19_2# comparator_equal_0/A3B3 0.08fF
C1214 GND comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.23fF
C1215 enable_2/enable 2_input_OR_0/w_30_15# 0.03fF
C1216 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C1217 VDD enable_2/2_input_AND_6/OUT 0.06fF
C1218 enable_1/2_input_AND_4/w_35_9# enable_1/2_input_AND_4/OUT 0.08fF
C1219 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1220 VDD adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# 0.03fF
C1221 VDD adder_subtractor_0/full_adder_1/2_input_OR_0/w_30_15# 0.03fF
C1222 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1223 and_block_0/2_input_AND_0/w_35_9# VDD 0.03fF
C1224 comparator_equal_0/4_input_AND_1/w_n22_4# comparator_equal_0/A2B2 0.07fF
C1225 comparator_equal_0/4_input_AND_0/w_n22_4# comparator_equal_0/4_input_AND_0/OUT 0.09fF
C1226 adder_subtractor_0/full_adder_3/2_input_AND_0/w_35_9# adder_subtractor_0/full_adder_3/2_input_AND_0/OUT 0.08fF
C1227 OUTPUT_ALU_ADDER_A3 adder_subtractor_0/B3_XOR 0.96fF
C1228 adder_subtractor_0/full_adder_2/2_input_OR_0/B adder_subtractor_0/full_adder_2/2_input_AND_0/w_35_9# 0.03fF
C1229 adder_subtractor_0/B1_XOR adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.12fF
C1230 and_block_0/2_input_AND_1/w_35_9# AND_OUTPUT_A1B1 0.04fF
C1231 GND comparator_equal_0/A3B3 0.83fF
C1232 GND enable_0/2_input_AND_2/OUT 0.04fF
C1233 VDD ADDER_SUB_C4 0.04fF
C1234 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# comparator_equal_0/A2B2 0.07fF
C1235 enable_0/2_input_AND_4/w_n12_9# INPUT_ALU_B0 0.07fF
C1236 comparator_equal_0/q1b_5_INPUT_AND_1/w_50_10# comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.07fF
C1237 comparator_equal_0/q1a_NOT_2/vdd comparator_equal_0/A2B2 0.11fF
C1238 VDD enable_1/2_input_AND_7/OUT 0.06fF
C1239 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_4/w_52_34# 0.09fF
C1240 GND adder_subtractor_0/full_adder_2/2_input_AND_0/OUT 0.04fF
C1241 VDD enable_2/2_input_AND_1/w_35_9# 0.03fF
C1242 enable_0/2_input_AND_4/OUT OUTPUT_ALU_ANDBLOCK_B0 0.05fF
C1243 comparator_equal_0/q1b_5_INPUT_AND_0/OUT comparator_equal_0/A2B2 0.17fF
C1244 VDD enable_1/2_input_AND_1/w_35_9# 0.03fF
C1245 INPUT_ALU_A3 decoder_0/A1_BAR 0.22fF
C1246 ADD_SUB_M ADDER_SUB_CFINAL 0.18fF
C1247 comparator_equal_0/A3NOT_B3 comparator_equal_0/2_input_AND_1/OUT 0.05fF
C1248 S0_S1_DECODER enable_0/2_input_AND_4/w_n12_9# 0.07fF
C1249 GND OUTPUT_ALU_ADDER_A1 1.22fF
C1250 OUTPUT_ALU_ANDBLOCK_A1 GND 0.32fF
C1251 comparator_equal_0/3_input_AND_1/w_n19_2# comparator_equal_0/A2NOT 0.08fF
C1252 VDD enable_2/2_input_AND_5/OUT 0.06fF
C1253 enable_1/2_input_AND_6/OUT OUTPUT_ALU_COMPARATOR_B2 0.05fF
C1254 enable_1/2_input_AND_5/w_35_9# OUTPUT_ALU_COMPARATOR_B1 0.03fF
C1255 VDD S0_DECODER 0.31fF
C1256 comparator_equal_0/B1_NOT comparator_equal_0/q1a_NOT_2/w_n12_4# 0.04fF
C1257 GND comparator_equal_0/A0NOT 0.27fF
C1258 VDD comparator_equal_0/q1a_NOT_6/w_n12_4# 0.05fF
C1259 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR 0.09fF
C1260 comparator_equal_0/A0B0 OUTPUT_ALU_COMPARATOR_A2 0.26fF
C1261 VDD comparator_equal_0/2_input_AND_1/w_35_9# 0.03fF
C1262 and_block_0/2_input_AND_3/w_35_9# and_block_0/2_input_AND_3/OUT 0.08fF
C1263 comparator_equal_0/B2_NOT comparator_equal_0/A3B3 0.50fF
C1264 ADDER_SUB_S1 ADDER_SUB_C1 0.15fF
C1265 adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.05fF
C1266 adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_2/2_input_OR_0/OUT 0.03fF
C1267 GND comparator_equal_0/A2NOT 0.47fF
C1268 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1269 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1270 VDD enable_0/2_input_AND_7/w_n12_9# 0.07fF
C1271 GND adder_subtractor_0/full_adder_2/2_input_OR_0/OUT 0.15fF
C1272 comparator_equal_0/A2_B2NOT_A3B3XNOR OUTPUT_ALU_COMPARATOR_B3 0.54fF
C1273 comparator_equal_0/XNOR_1/OUT comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C1274 GND OUTPUT_ALU_ANDBLOCK_B2 0.40fF
C1275 comparator_equal_0/4_input_AND_1/w_n22_4# comparator_equal_0/4_input_AND_1/OUT 0.09fF
C1276 VDD S0BAR_S1_DECODER 0.69fF
C1277 INPUT_ALU_B2 enable_2/2_input_AND_6/OUT 0.02fF
C1278 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.08fF
C1279 INPUT_ALU_A2 decoder_0/A1_BAR 0.28fF
C1280 comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/q1a_NOT_2/vdd 0.21fF
C1281 GND comparator_equal_0/B0_NOT 0.10fF
C1282 GND adder_subtractor_0/full_adder_1/2_input_OR_0/A 0.44fF
C1283 VDD enable_2/2_input_AND_4/OUT 0.06fF
C1284 decoder_0/2_input_AND_1/OUT decoder_0/2_input_AND_1/w_n12_9# 0.03fF
C1285 enable_1/2_input_AND_3/w_35_9# enable_1/2_input_AND_3/OUT 0.08fF
C1286 VDD adder_subtractor_0/q1d_2_INPUT_XOR_3/w_12_2# 0.03fF
C1287 OUTPUT_ALU_ANDBLOCK_A0 GND 0.10fF
C1288 comparator_equal_0/4_input_AND_0/w_n22_4# comparator_equal_0/A3B3 0.07fF
C1289 comparator_equal_0/A3NOT_B3 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C1290 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 2.05fF
C1291 VDD comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C1292 comparator_equal_0/A1B1 OUTPUT_ALU_COMPARATOR_A2 0.27fF
C1293 adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_0/2_input_AND_1/OUT 0.03fF
C1294 VDD adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR 0.03fF
C1295 adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# ADDER_SUB_C2 0.07fF
C1296 enable_2/enable INPUT_ALU_A1 0.66fF
C1297 AND_OUTPUT_A3B3 VDD 0.02fF
C1298 comparator_equal_0/4_input_AND_0/OUT comparator_equal_0/A2B2 0.09fF
C1299 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.17fF
C1300 adder_subtractor_0/full_adder_3/2_input_OR_0/A adder_subtractor_0/full_adder_3/2_input_OR_0/B 0.45fF
C1301 adder_subtractor_0/full_adder_3/2_input_OR_0/w_30_15# adder_subtractor_0/full_adder_3/2_input_OR_0/OUT 0.06fF
C1302 adder_subtractor_0/full_adder_1/2_input_OR_0/B adder_subtractor_0/full_adder_1/2_input_OR_0/OUT 0.20fF
C1303 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A2_B2NOT_A3B3XNOR 0.35fF
C1304 VDD comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1305 GND 2_input_AND_0/OUT 0.04fF
C1306 VDD comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# 0.11fF
C1307 enable_2/2_input_AND_1/w_35_9# enable_2/2_input_AND_1/OUT 0.08fF
C1308 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1309 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C1310 ADDER_SUB_S0 GND 0.33fF
C1311 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_0/AXORB 0.19fF
C1312 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_53_n17# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C1313 and_block_0/2_input_AND_0/w_35_9# AND_OUTPUT_A0B0 0.03fF
C1314 GND OUTPUT_ALU_ANDBLOCK_B1 0.34fF
C1315 VDD adder_subtractor_0/full_adder_2/2_input_AND_1/w_35_9# 0.03fF
C1316 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_53_n17# 0.03fF
C1317 ADD_SUB_M VDD 2.15fF
C1318 VDD decoder_0/2_input_AND_0/w_n12_9# 0.06fF
C1319 enable_1/2_input_AND_4/OUT OUTPUT_ALU_COMPARATOR_B0 0.05fF
C1320 enable_0/2_input_AND_3/w_35_9# enable_0/2_input_AND_3/OUT 0.08fF
C1321 2_input_OR_0/a_n7_22# INPUT_ALU_B1 0.00fF
C1322 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_ADDER_A3 0.03fF
C1323 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR VDD 0.03fF
C1324 VDD enable_2/2_input_AND_3/OUT 0.06fF
C1325 GND OUTPUT_ALU_COMPARATOR_B3 1.55fF
C1326 GND adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR 0.04fF
C1327 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.03fF
C1328 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_S0 0.03fF
C1329 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 comparator_equal_0/A3B3 0.30fF
C1330 OUTPUT_ALU_ADDER_B0 enable_2/2_input_AND_4/OUT 0.05fF
C1331 enable_1/2_input_AND_7/w_n12_9# INPUT_ALU_B3 0.07fF
C1332 COMPARATOR_A_EQUAL_B_FINAL 2_input_AND_0/w_35_9# 0.03fF
C1333 VDD adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_n34_1# 0.03fF
C1334 INPUT_ALU_A3 decoder_0/2_input_AND_0/a_4_n21# 0.00fF
C1335 S0_DECODER S0BAR_S1BAR_DECODER 0.12fF
C1336 S0BAR_S1_DECODER enable_1/2_input_AND_6/OUT 0.12fF
C1337 adder_subtractor_0/B0_XOR ADD_SUB_M 0.18fF
C1338 adder_subtractor_0/full_adder_1/2_input_AND_1/w_35_9# adder_subtractor_0/full_adder_1/2_input_AND_1/OUT 0.08fF
C1339 ADDER_SUB_C1 adder_subtractor_0/full_adder_1/AXORB 0.93fF
C1340 decoder_0/2_input_AND_1/OUT S0_DECODER 0.12fF
C1341 OUTPUT_ALU_ADDER_B2 adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 1.31fF
C1342 adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# adder_subtractor_0/full_adder_3/AXORB 0.07fF
C1343 and_block_0/2_input_AND_2/w_35_9# and_block_0/2_input_AND_2/OUT 0.08fF
C1344 enable_2/2_input_AND_1/w_n12_9# enable_2/enable 0.07fF
C1345 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/full_adder_2/AXORB 0.03fF
C1346 AND_OUTPUT_A2B2 VDD 0.02fF
C1347 VDD comparator_equal_0/B3_NOT 0.10fF
C1348 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_52_34# ADDER_SUB_C3 0.09fF
C1349 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C1350 comparator_equal_0/3_input_AND_0/w_n19_2# comparator_equal_0/B2_NOT 0.08fF
C1351 S0BAR_S1_DECODER INPUT_ALU_B2 0.55fF
C1352 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR OUTPUT_ALU_ADDER_A0 0.11fF
C1353 S0BAR_S1_DECODER enable_1/2_input_AND_1/w_n12_9# 0.07fF
C1354 GND adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR 0.04fF
C1355 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/A2B2 0.34fF
C1356 GND OUTPUT_ALU_ANDBLOCK_B0 0.16fF
C1357 OUTPUT_ALU_ADDER_A1 comparator_equal_0/A1NOTB1_A2XNORB2_A3XNORB3 0.20fF
C1358 comparator_equal_0/XNOR_3/OUT comparator_equal_0/XNOR_3/w_181_105# 0.13fF
C1359 adder_subtractor_0/B0_XOR VDD 0.37fF
C1360 comparator_equal_0/2_input_AND_0/w_n12_9# comparator_equal_0/2_input_AND_0/OUT 0.03fF
C1361 VDD adder_subtractor_0/full_adder_2/2_input_AND_0/w_35_9# 0.03fF
C1362 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# 0.09fF
C1363 VDD comparator_equal_0/4_input_AND_2/OUT 0.21fF
C1364 comparator_equal_0/3_input_AND_0/OUT OUTPUT_ALU_COMPARATOR_A2 0.13fF
C1365 OUTPUT_ALU_COMPARATOR_B0 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# 0.08fF
C1366 GND OUTPUT_ALU_COMPARATOR_A3 1.02fF
C1367 ADD_SUB_M OUTPUT_ALU_ADDER_B0 0.42fF
C1368 adder_subtractor_0/B2_XOR adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.19fF
C1369 decoder_0/A0_BAR S0_DECODER 0.04fF
C1370 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_0/AXORB 0.08fF
C1371 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.10fF
C1372 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/XNOR_3/OUT 0.15fF
C1373 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_12_2# adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C1374 VDD enable_2/2_input_AND_2/OUT 0.06fF
C1375 OUTPUT_ALU_COMPARATOR_A0 enable_1/2_input_AND_0/w_35_9# 0.13fF
C1376 comparator_equal_0/4_input_AND_2/w_n22_4# comparator_equal_0/A1NOT 0.07fF
C1377 comparator_equal_0/A2NOT_B2_A3B3XNOR comparator_equal_0/3_input_AND_1/OUT 0.05fF
C1378 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR comparator_equal_0/q1c_4_INPUT_OR_0/OUT 0.78fF
C1379 comparator_equal_0/A3B3 comparator_equal_0/A2B2 5.18fF
C1380 INPUT_ALU_A1 S1_DECODER 0.06fF
C1381 GND comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.23fF
C1382 S0BAR_S1_DECODER enable_1/2_input_AND_5/OUT 0.12fF
C1383 adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# adder_subtractor_0/full_adder_0/2_input_AND_0/OUT 0.03fF
C1384 VDD OUTPUT_ALU_ADDER_B0 1.53fF
C1385 OUTPUT_ALU_ADDER_A0 enable_2/2_input_AND_0/w_35_9# 0.14fF
C1386 adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# OUTPUT_ALU_ADDER_A2 0.07fF
C1387 OUTPUT_ALU_ADDER_A1 adder_subtractor_0/full_adder_1/AXORB 0.15fF
C1388 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_53_n17# adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR 0.03fF
C1389 INPUT_ALU_A1 decoder_0/2_input_AND_2/OUT 0.05fF
C1390 VDD enable_0/2_input_AND_1/OUT 0.06fF
C1391 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_52_34# adder_subtractor_0/B2_XOR 0.03fF
C1392 AND_OUTPUT_A1B1 VDD 0.02fF
C1393 decoder_0/2_input_AND_0/OUT decoder_0/2_input_AND_0/w_n12_9# 0.03fF
C1394 ADD_SUB_M INPUT_ALU_B2 0.51fF
C1395 GND ADDER_SUB_C2 0.80fF
C1396 GND adder_subtractor_0/full_adder_0/AXORB 0.33fF
C1397 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C1398 comparator_equal_0/2_input_AND_1/w_35_9# comparator_equal_0/2_input_AND_1/OUT 0.08fF
C1399 OUTPUT_ALU_COMPARATOR_B3 comparator_equal_0/2_input_AND_1/w_n12_9# 0.07fF
C1400 S0BAR_S1_DECODER INPUT_ALU_B1 0.66fF
C1401 GND INPUT_ALU_A1 2.74fF
C1402 VDD comparator_equal_0/3_input_AND_1/w_34_3# 0.03fF
C1403 ADDER_SUB_S3 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR 0.19fF
C1404 VDD enable_1/2_input_AND_6/OUT 0.06fF
C1405 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# comparator_equal_0/A3B3 0.09fF
C1406 GND OUTPUT_ALU_ANDBLOCK_B3 0.32fF
C1407 VDD adder_subtractor_0/full_adder_2/2_input_OR_0/w_30_15# 0.03fF
C1408 adder_subtractor_0/full_adder_0/2_input_OR_0/A VDD 0.18fF
C1409 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/XNOR_3/OUT 0.18fF
C1410 ADD_SUB_M S0BAR_S1BAR_DECODER 0.67fF
C1411 VDD decoder_0/2_input_AND_0/OUT 0.06fF
C1412 adder_subtractor_0/B0_XOR OUTPUT_ALU_ADDER_B0 0.21fF
C1413 ADD_SUB_M decoder_0/2_input_AND_1/OUT 0.05fF
C1414 VDD enable_2/2_input_AND_0/OUT 0.06fF
C1415 enable_2/enable 2_input_OR_0/OUT 0.05fF
C1416 adder_subtractor_0/B2_XOR adder_subtractor_0/B3_XOR 0.15fF
C1417 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT ADDER_SUB_C3 0.05fF
C1418 OUTPUT_ALU_COMPARATOR_B0 OUTPUT_ALU_COMPARATOR_B1 0.14fF
C1419 comparator_equal_0/q1b_5_INPUT_AND_1/OUT comparator_equal_0/A3B3 0.05fF
C1420 comparator_equal_0/A0NOT comparator_equal_0/A2B2 0.08fF
C1421 VDD INPUT_ALU_B2 0.18fF
C1422 OUTPUT_ALU_COMPARATOR_A0 OUTPUT_ALU_COMPARATOR_B1 0.47fF
C1423 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_53_n17# ADDER_SUB_S3 0.04fF
C1424 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/4_input_AND_1/OUT 0.14fF
C1425 VDD enable_1/2_input_AND_1/w_n12_9# 0.06fF
C1426 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_52_34# adder_subtractor_0/full_adder_0/AXORB 0.03fF
C1427 VDD enable_2/2_input_AND_1/OUT 0.06fF
C1428 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR OUTPUT_ALU_ADDER_B1 0.03fF
C1429 GND adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR 0.25fF
C1430 OUTPUT_ALU_COMPARATOR_B2 OUTPUT_ALU_COMPARATOR_B1 0.08fF
C1431 GND comparator_equal_0/A0B0 1.64fF
C1432 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_53_n17# ADDER_SUB_S0 0.04fF
C1433 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_12_2# adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C1434 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C1435 VDD comparator_equal_0/q1a_NOT_5/in 0.44fF
C1436 S0BAR_S1_DECODER enable_1/2_input_AND_4/OUT 0.12fF
C1437 VDD S0BAR_S1BAR_DECODER 0.02fF
C1438 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_2/AXORB 0.08fF
C1439 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_12_2# ADDER_SUB_C2 0.08fF
C1440 adder_subtractor_0/full_adder_1/2_input_AND_0/w_35_9# adder_subtractor_0/full_adder_1/2_input_AND_0/OUT 0.08fF
C1441 OUTPUT_ALU_ADDER_A1 adder_subtractor_0/B1_XOR 0.90fF
C1442 adder_subtractor_0/full_adder_0/2_input_OR_0/B adder_subtractor_0/full_adder_0/2_input_AND_0/w_35_9# 0.03fF
C1443 adder_subtractor_0/full_adder_3/2_input_OR_0/A adder_subtractor_0/full_adder_3/2_input_AND_1/w_35_9# 0.03fF
C1444 adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# adder_subtractor_0/B3_XOR 0.07fF
C1445 and_block_0/2_input_AND_1/w_35_9# and_block_0/2_input_AND_1/OUT 0.08fF
C1446 VDD decoder_0/2_input_AND_1/OUT 0.06fF
C1447 GND comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.14fF
C1448 S0BAR_S1_DECODER enable_1/2_input_AND_0/w_n12_9# 0.07fF
C1449 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# comparator_equal_0/A0NOT 0.07fF
C1450 comparator_equal_0/q1b_5_INPUT_AND_0/w_50_10# comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 0.04fF
C1451 S0BAR_S1_DECODER COMPARATOR_OUT_A_EQUAL_B 0.79fF
C1452 AND_OUTPUT_A0B0 VDD 0.02fF
C1453 ADD_SUB_M INPUT_ALU_B1 0.87fF
C1454 comparator_equal_0/B1_NOT OUTPUT_ALU_COMPARATOR_B1 0.04fF
C1455 comparator_equal_0/4_input_AND_1/OUT comparator_equal_0/A3B3 0.15fF
C1456 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR ADDER_SUB_C2 0.51fF
C1457 GND OUTPUT_ALU_ADDER_A2 1.29fF
C1458 GND OUTPUT_ALU_ADDER_A0 1.91fF
C1459 decoder_0/A0_BAR decoder_0/2_input_AND_0/w_n12_9# 0.07fF
C1460 S0BAR_S1_DECODER INPUT_ALU_B0 0.66fF
C1461 comparator_equal_0/q1a_NOT_5/in comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR 0.40fF
C1462 VDD enable_2/2_input_AND_7/OUT 0.06fF
C1463 VDD comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C1464 VDD enable_1/2_input_AND_5/OUT 0.06fF
C1465 enable_0/2_input_AND_7/w_n12_9# S0_S1_DECODER 0.07fF
C1466 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/q1d_2_INPUT_XOR_1/w_n34_1# 0.03fF
C1467 comparator_equal_0/A0NOT comparator_equal_0/q1b_5_INPUT_AND_1/OUT 0.13fF
C1468 comparator_equal_0/B0_NOT comparator_equal_0/A2B2 0.08fF
C1469 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_12_2# VDD 0.03fF
C1470 VDD comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1471 INPUT_ALU_A3 S0_DECODER 0.17fF
C1472 VDD decoder_0/A0_BAR 0.32fF
C1473 VDD INPUT_ALU_B1 0.30fF
C1474 OUTPUT_ALU_ADDER_B2 INPUT_ALU_B3 0.05fF
C1475 OUTPUT_ALU_COMPARATOR_A1 comparator_equal_0/q1a_NOT_7/w_n12_4# 0.12fF
C1476 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_n34_1# adder_subtractor_0/B3_XOR 0.08fF
C1477 GND comparator_equal_0/A1B1 1.87fF
C1478 GND OUTPUT_ALU_ADDER_B1 1.48fF
C1479 comparator_equal_0/A2NOT comparator_equal_0/3_input_AND_1/OUT 0.13fF
C1480 S0BAR_S1_DECODER enable_1/2_input_AND_3/OUT 0.12fF
C1481 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# 0.07fF
C1482 adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_0/2_input_OR_0/OUT 0.03fF
C1483 comparator_equal_0/A2_B2NOT_A3B3XNOR comparator_equal_0/3_input_AND_0/OUT 0.05fF
C1484 adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_2/2_input_OR_0/A 0.07fF
C1485 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# comparator_equal_0/XNOR_1/OUT 0.03fF
C1486 VDD adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR 0.03fF
C1487 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_n34_1# adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1488 VDD comparator_equal_0/2_input_AND_1/OUT 0.06fF
C1489 VDD enable_0/2_input_AND_0/w_35_9# 0.03fF
C1490 and_block_0/2_input_AND_3/OUT AND_OUTPUT_A3B3 0.05fF
C1491 ADD_SUB_M INPUT_ALU_B0 0.29fF
C1492 OUTPUT_ALU_COMPARATOR_A0 comparator_equal_0/q1b_5_INPUT_AND_0/OUT 0.13fF
C1493 GND adder_subtractor_0/full_adder_2/2_input_OR_0/A 0.44fF
C1494 adder_subtractor_0/full_adder_0/2_input_OR_0/B GND 0.16fF
C1495 S0BAR_S1_DECODER INPUT_ALU_A3 0.64fF
C1496 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# 0.03fF
C1497 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR adder_subtractor_0/full_adder_3/AXORB 0.24fF
C1498 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_53_n17# adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR 0.03fF
C1499 GND enable_0/2_input_AND_6/OUT 0.04fF
C1500 decoder_0/q1a_NOT_1/w_n12_4# S1_DECODER 0.07fF
C1501 enable_0/2_input_AND_7/OUT OUTPUT_ALU_ANDBLOCK_B3 0.05fF
C1502 comparator_equal_0/4_input_AND_1/w_n22_4# comparator_equal_0/B1_NOT 0.08fF
C1503 VDD enable_1/2_input_AND_4/OUT 0.06fF
C1504 VDD comparator_equal_0/4_input_AND_0/w_40_5# 0.03fF
C1505 enable_2/2_input_AND_6/w_n12_9# enable_2/2_input_AND_6/OUT 0.03fF
C1506 comparator_equal_0/A2B2 OUTPUT_ALU_COMPARATOR_B3 0.73fF
C1507 GND enable_1/2_input_AND_1/OUT 0.04fF
C1508 VDD enable_1/2_input_AND_0/w_n12_9# 0.06fF
C1509 comparator_equal_0/B1_NOT comparator_equal_0/q1a_NOT_2/vdd 0.10fF
C1510 comparator_equal_0/4_input_AND_0/w_n22_4# comparator_equal_0/A0B0 0.07fF
C1511 VDD COMPARATOR_OUT_A_EQUAL_B 0.22fF
C1512 enable_0/2_input_AND_1/w_n12_9# INPUT_ALU_A1 0.07fF
C1513 INPUT_ALU_A2 S0_DECODER 0.17fF
C1514 decoder_0/2_input_AND_0/OUT S0BAR_S1BAR_DECODER 0.05fF
C1515 VDD INPUT_ALU_B0 0.37fF
C1516 VDD adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# 0.24fF
C1517 OUTPUT_ALU_ADDER_B0 INPUT_ALU_B1 0.05fF
C1518 comparator_equal_0/A3NOT_B3 comparator_equal_0/A2NOT_B2_A3B3XNOR 2.38fF
C1519 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C1520 OUTPUT_ALU_ADDER_B1 enable_2/2_input_AND_5/w_35_9# 0.03fF
C1521 enable_0/2_input_AND_3/w_n12_9# enable_0/2_input_AND_3/OUT 0.03fF
C1522 GND 2_input_OR_0/OUT 0.15fF
C1523 adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# ADD_SUB_M 0.07fF
C1524 VDD enable_0/2_input_AND_0/w_n12_9# 0.06fF
C1525 S0BAR_S1_DECODER enable_1/2_input_AND_2/OUT 0.12fF
C1526 and_block_0/2_input_AND_3/OUT VDD 0.06fF
C1527 comparator_equal_0/q1c_4_INPUT_OR_1/w_41_n9# COMPARATOR_OUT_A_LESSTHAN_B 0.05fF
C1528 comparator_equal_0/A3NOT_B3 comparator_equal_0/q1c_4_INPUT_OR_1/OUT 0.09fF
C1529 adder_subtractor_0/full_adder_1/2_input_OR_0/A adder_subtractor_0/full_adder_1/2_input_OR_0/B 0.45fF
C1530 adder_subtractor_0/full_adder_1/2_input_OR_0/w_30_15# adder_subtractor_0/full_adder_1/2_input_OR_0/OUT 0.06fF
C1531 adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# adder_subtractor_0/full_adder_3/2_input_OR_0/B 0.07fF
C1532 INPUT_ALU_B3 OUTPUT_ALU_COMPARATOR_B2 0.07fF
C1533 VDD S0_S1_DECODER 0.02fF
C1534 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/2_input_AND_0/OUT 0.12fF
C1535 adder_subtractor_0/full_adder_2/AXORB adder_subtractor_0/full_adder_2/2_input_AND_1/OUT 0.12fF
C1536 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/q1a_NOT_1/w_n12_4# 0.10fF
C1537 ADD_SUB_M INPUT_ALU_A3 0.24fF
C1538 GND enable_1/2_input_AND_0/OUT 0.04fF
C1539 OUTPUT_ALU_COMPARATOR_A3 comparator_equal_0/A2B2 0.16fF
C1540 OUTPUT_ALU_COMPARATOR_B2 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C1541 VDD comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C1542 S0BAR_S1_DECODER INPUT_ALU_A2 0.71fF
C1543 and_block_0/2_input_AND_0/w_35_9# and_block_0/2_input_AND_0/OUT 0.08fF
C1544 INPUT_ALU_A3 decoder_0/2_input_AND_0/w_n12_9# 0.02fF
C1545 decoder_0/A0_BAR decoder_0/2_input_AND_0/OUT 0.12fF
C1546 GND enable_0/2_input_AND_5/OUT 0.04fF
C1547 adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# VDD 0.06fF
C1548 GND comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.23fF
C1549 VDD enable_1/2_input_AND_3/OUT 0.06fF
C1550 GND comparator_equal_0/3_input_AND_0/OUT 0.09fF
C1551 VDD comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.07fF
C1552 INPUT_ALU_B1 INPUT_ALU_B2 0.85fF
C1553 GND OUTPUT_ALU_COMPARATOR_A2 1.00fF
C1554 OUTPUT_ALU_ADDER_A2 OUTPUT_ALU_ADDER_B3 0.38fF
C1555 ADD_SUB_M adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR 0.08fF
C1556 comparator_equal_0/A1B1 comparator_equal_0/4_input_AND_0/w_n22_4# 0.08fF
C1557 VDD enable_1/2_input_AND_0/w_35_9# 0.03fF
C1558 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR VDD 0.03fF
C1559 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR OUTPUT_ALU_COMPARATOR_B1 0.03fF
C1560 VDD INPUT_ALU_A3 0.69fF
C1561 INPUT_ALU_B1 S0BAR_S1BAR_DECODER 0.44fF
C1562 S0_DECODER decoder_0/q1a_NOT_0/w_n12_4# 0.07fF
C1563 COMPARATOR_A_EQUAL_B_FINAL 2_input_AND_0/OUT 0.05fF
C1564 GND adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR 0.04fF
C1565 GND adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR 0.27fF
C1566 decoder_0/q1a_NOT_1/w_n12_4# Gnd 0.50fF
C1567 decoder_0/q1a_NOT_0/w_n12_4# Gnd 0.50fF
C1568 decoder_0/2_input_AND_3/OUT Gnd 0.38fF
C1569 decoder_0/2_input_AND_3/w_35_9# Gnd 0.56fF
C1570 decoder_0/2_input_AND_3/w_n12_9# Gnd 0.72fF
C1571 decoder_0/2_input_AND_2/OUT Gnd 0.38fF
C1572 decoder_0/2_input_AND_2/w_35_9# Gnd 0.56fF
C1573 decoder_0/2_input_AND_2/w_n12_9# Gnd 0.72fF
C1574 decoder_0/2_input_AND_1/OUT Gnd 0.38fF
C1575 S0_DECODER Gnd 2.34fF
C1576 decoder_0/A1_BAR Gnd 0.50fF
C1577 decoder_0/2_input_AND_1/w_35_9# Gnd 0.56fF
C1578 decoder_0/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1579 S0BAR_S1BAR_DECODER Gnd 1.54fF
C1580 decoder_0/2_input_AND_0/OUT Gnd 0.38fF
C1581 decoder_0/A0_BAR Gnd 1.04fF
C1582 decoder_0/2_input_AND_0/w_35_9# Gnd 0.56fF
C1583 decoder_0/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1584 comparator_equal_0/q1a_NOT_2/w_n12_4# Gnd 0.50fF
C1585 comparator_equal_0/q1a_NOT_1/w_n12_4# Gnd 0.50fF
C1586 comparator_equal_0/q1a_NOT_0/w_n12_4# Gnd 0.50fF
C1587 comparator_equal_0/XNOR_3/w_181_105# Gnd 2.32fF
C1588 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1589 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1590 comparator_equal_0/XNOR_3/OUT Gnd 1.20fF
C1591 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1592 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1593 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1594 comparator_equal_0/XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1595 comparator_equal_0/2_input_AND_1/OUT Gnd 0.38fF
C1596 comparator_equal_0/q1a_NOT_4/out Gnd 0.58fF
C1597 OUTPUT_ALU_COMPARATOR_B3 Gnd 2.65fF
C1598 comparator_equal_0/2_input_AND_1/w_35_9# Gnd 0.56fF
C1599 comparator_equal_0/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1600 comparator_equal_0/XNOR_2/w_181_105# Gnd 2.32fF
C1601 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1602 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1603 comparator_equal_0/XNOR_2/OUT Gnd 1.20fF
C1604 OUTPUT_ALU_COMPARATOR_A2 Gnd 8.37fF
C1605 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1606 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1607 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1608 comparator_equal_0/XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1609 comparator_equal_0/4_input_AND_2/OUT Gnd 0.72fF
C1610 comparator_equal_0/A1NOT Gnd 0.93fF
C1611 OUTPUT_ALU_COMPARATOR_B1 Gnd 1.94fF
C1612 comparator_equal_0/A2B2 Gnd 2.49fF
C1613 comparator_equal_0/A3B3 Gnd 3.25fF
C1614 comparator_equal_0/4_input_AND_2/w_40_5# Gnd 0.51fF
C1615 comparator_equal_0/4_input_AND_2/w_n22_4# Gnd 0.99fF
C1616 comparator_equal_0/3_input_AND_1/OUT Gnd 0.51fF
C1617 comparator_equal_0/A2NOT Gnd 0.94fF
C1618 OUTPUT_ALU_COMPARATOR_B2 Gnd 1.83fF
C1619 comparator_equal_0/3_input_AND_1/w_34_3# Gnd 0.48fF
C1620 comparator_equal_0/3_input_AND_1/w_n19_2# Gnd 0.83fF
C1621 comparator_equal_0/2_input_AND_0/OUT Gnd 0.38fF
C1622 comparator_equal_0/B3_NOT Gnd 0.41fF
C1623 comparator_equal_0/2_input_AND_0/w_35_9# Gnd 0.56fF
C1624 comparator_equal_0/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1625 comparator_equal_0/A0B0 Gnd 1.50fF
C1626 comparator_equal_0/XNOR_0/w_181_105# Gnd 2.32fF
C1627 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1628 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1629 comparator_equal_0/XNOR_0/OUT Gnd 1.20fF
C1630 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1631 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1632 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1633 comparator_equal_0/XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1634 comparator_equal_0/XNOR_1/w_181_105# Gnd 2.32fF
C1635 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1636 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1637 comparator_equal_0/XNOR_1/OUT Gnd 1.20fF
C1638 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1639 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1640 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1641 comparator_equal_0/XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1642 comparator_equal_0/q1a_NOT_2/vdd Gnd 0.59fF
C1643 comparator_equal_0/4_input_AND_1/OUT Gnd 0.72fF
C1644 comparator_equal_0/B1_NOT Gnd 0.67fF
C1645 comparator_equal_0/4_input_AND_1/w_40_5# Gnd 0.51fF
C1646 comparator_equal_0/4_input_AND_1/w_n22_4# Gnd 0.99fF
C1647 comparator_equal_0/3_input_AND_0/OUT Gnd 0.51fF
C1648 comparator_equal_0/B2_NOT Gnd 0.41fF
C1649 comparator_equal_0/3_input_AND_0/w_34_3# Gnd 0.48fF
C1650 comparator_equal_0/3_input_AND_0/w_n19_2# Gnd 0.83fF
C1651 COMPARATOR_OUT_A_EQUAL_B Gnd 0.57fF
C1652 comparator_equal_0/4_input_AND_0/OUT Gnd 0.72fF
C1653 comparator_equal_0/4_input_AND_0/w_40_5# Gnd 0.51fF
C1654 comparator_equal_0/4_input_AND_0/w_n22_4# Gnd 0.99fF
C1655 COMPARATOR_OUT_A_LESSTHAN_B Gnd 0.37fF
C1656 comparator_equal_0/q1c_4_INPUT_OR_1/OUT Gnd 0.92fF
C1657 comparator_equal_0/A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 Gnd 7.27fF
C1658 comparator_equal_0/A2NOT_B2_A3B3XNOR Gnd 4.26fF
C1659 comparator_equal_0/A3NOT_B3 Gnd 4.30fF
C1660 comparator_equal_0/q1c_4_INPUT_OR_1/w_41_n9# Gnd 1.25fF
C1661 comparator_equal_0/q1c_4_INPUT_OR_1/w_n38_n10# Gnd 1.97fF
C1662 COMPARATOR_OUT_A_GREATERTHAN_B Gnd 0.53fF
C1663 comparator_equal_0/q1c_4_INPUT_OR_0/OUT Gnd 0.92fF
C1664 comparator_equal_0/A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR Gnd 13.09fF
C1665 comparator_equal_0/A1_B1NOT_A3B3XNOR_A2B2XOR Gnd 16.15fF
C1666 comparator_equal_0/A2_B2NOT_A3B3XNOR Gnd 7.25fF
C1667 comparator_equal_0/A3_B3NOT Gnd 1.55fF
C1668 comparator_equal_0/q1c_4_INPUT_OR_0/w_41_n9# Gnd 1.25fF
C1669 comparator_equal_0/q1c_4_INPUT_OR_0/w_n38_n10# Gnd 1.97fF
C1670 comparator_equal_0/q1b_5_INPUT_AND_1/OUT Gnd 0.31fF
C1671 comparator_equal_0/A0NOT Gnd 0.71fF
C1672 comparator_equal_0/A1B1 Gnd 1.91fF
C1673 comparator_equal_0/q1b_5_INPUT_AND_1/w_50_10# Gnd 0.06fF
C1674 comparator_equal_0/q1b_5_INPUT_AND_1/w_n24_8# Gnd 1.35fF
C1675 comparator_equal_0/q1b_5_INPUT_AND_0/OUT Gnd 0.31fF
C1676 comparator_equal_0/B0_NOT Gnd 0.42fF
C1677 comparator_equal_0/q1b_5_INPUT_AND_0/w_50_10# Gnd 0.06fF
C1678 comparator_equal_0/q1b_5_INPUT_AND_0/w_n24_8# Gnd 1.35fF
C1679 OUTPUT_ALU_COMPARATOR_A1 Gnd 10.85fF
C1680 comparator_equal_0/q1a_NOT_7/w_n12_4# Gnd 0.50fF
C1681 OUTPUT_ALU_COMPARATOR_A0 Gnd 15.75fF
C1682 comparator_equal_0/q1a_NOT_6/w_n12_4# Gnd 0.50fF
C1683 comparator_equal_0/q1a_NOT_5/in Gnd 0.49fF
C1684 comparator_equal_0/q1a_NOT_5/w_n12_4# Gnd 0.50fF
C1685 OUTPUT_ALU_COMPARATOR_A3 Gnd 4.53fF
C1686 comparator_equal_0/q1a_NOT_4/w_n12_4# Gnd 0.50fF
C1687 comparator_equal_0/q1a_NOT_3/w_n12_4# Gnd 0.50fF
C1688 COMPARATOR_A_EQUAL_B_FINAL Gnd 0.14fF
C1689 2_input_AND_0/OUT Gnd 0.38fF
C1690 2_input_AND_0/w_35_9# Gnd 0.56fF
C1691 2_input_AND_0/w_n12_9# Gnd 0.72fF
C1692 enable_2/2_input_AND_6/OUT Gnd 0.38fF
C1693 INPUT_ALU_B2 Gnd 1.49fF
C1694 enable_2/2_input_AND_6/w_35_9# Gnd 0.56fF
C1695 enable_2/2_input_AND_6/w_n12_9# Gnd 0.72fF
C1696 enable_2/2_input_AND_5/OUT Gnd 0.38fF
C1697 INPUT_ALU_B1 Gnd 1.31fF
C1698 enable_2/2_input_AND_5/w_35_9# Gnd 0.56fF
C1699 enable_2/2_input_AND_5/w_n12_9# Gnd 0.72fF
C1700 enable_2/2_input_AND_4/OUT Gnd 0.38fF
C1701 INPUT_ALU_B0 Gnd 1.35fF
C1702 enable_2/2_input_AND_4/w_35_9# Gnd 0.56fF
C1703 enable_2/2_input_AND_4/w_n12_9# Gnd 0.72fF
C1704 enable_2/2_input_AND_3/OUT Gnd 0.38fF
C1705 INPUT_ALU_A3 Gnd 30.86fF
C1706 enable_2/2_input_AND_3/w_35_9# Gnd 0.56fF
C1707 enable_2/2_input_AND_3/w_n12_9# Gnd 0.72fF
C1708 enable_2/2_input_AND_2/OUT Gnd 0.38fF
C1709 INPUT_ALU_A2 Gnd 36.52fF
C1710 enable_2/2_input_AND_2/w_35_9# Gnd 0.56fF
C1711 enable_2/2_input_AND_2/w_n12_9# Gnd 0.72fF
C1712 enable_2/2_input_AND_1/OUT Gnd 0.38fF
C1713 INPUT_ALU_A1 Gnd 22.06fF
C1714 enable_2/2_input_AND_1/w_35_9# Gnd 0.56fF
C1715 enable_2/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1716 enable_2/2_input_AND_0/OUT Gnd 0.38fF
C1717 enable_2/enable Gnd 2.77fF
C1718 INPUT_ALU_A0 Gnd 31.80fF
C1719 enable_2/2_input_AND_0/w_35_9# Gnd 0.56fF
C1720 enable_2/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1721 enable_2/2_input_AND_7/OUT Gnd 0.38fF
C1722 INPUT_ALU_B3 Gnd 1.61fF
C1723 enable_2/2_input_AND_7/w_35_9# Gnd 0.56fF
C1724 enable_2/2_input_AND_7/w_n12_9# Gnd 0.72fF
C1725 2_input_OR_0/OUT Gnd 0.41fF
C1726 2_input_OR_0/w_30_15# Gnd 0.60fF
C1727 2_input_OR_0/w_n23_15# Gnd 0.73fF
C1728 enable_1/2_input_AND_6/OUT Gnd 0.38fF
C1729 enable_1/2_input_AND_6/w_35_9# Gnd 0.56fF
C1730 enable_1/2_input_AND_6/w_n12_9# Gnd 0.72fF
C1731 enable_1/2_input_AND_5/OUT Gnd 0.38fF
C1732 enable_1/2_input_AND_5/w_35_9# Gnd 0.56fF
C1733 enable_1/2_input_AND_5/w_n12_9# Gnd 0.72fF
C1734 enable_1/2_input_AND_4/OUT Gnd 0.38fF
C1735 enable_1/2_input_AND_4/w_35_9# Gnd 0.56fF
C1736 enable_1/2_input_AND_4/w_n12_9# Gnd 0.72fF
C1737 enable_1/2_input_AND_3/OUT Gnd 0.38fF
C1738 enable_1/2_input_AND_3/w_35_9# Gnd 0.56fF
C1739 enable_1/2_input_AND_3/w_n12_9# Gnd 0.72fF
C1740 enable_1/2_input_AND_2/OUT Gnd 0.38fF
C1741 enable_1/2_input_AND_2/w_35_9# Gnd 0.56fF
C1742 enable_1/2_input_AND_2/w_n12_9# Gnd 0.72fF
C1743 enable_1/2_input_AND_1/OUT Gnd 0.38fF
C1744 enable_1/2_input_AND_1/w_35_9# Gnd 0.56fF
C1745 enable_1/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1746 enable_1/2_input_AND_0/OUT Gnd 0.38fF
C1747 enable_1/2_input_AND_0/w_35_9# Gnd 0.56fF
C1748 enable_1/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1749 enable_1/2_input_AND_7/OUT Gnd 0.38fF
C1750 enable_1/2_input_AND_7/w_35_9# Gnd 0.56fF
C1751 enable_1/2_input_AND_7/w_n12_9# Gnd 0.72fF
C1752 OUTPUT_ALU_ANDBLOCK_B2 Gnd 0.70fF
C1753 enable_0/2_input_AND_6/OUT Gnd 0.38fF
C1754 enable_0/2_input_AND_6/w_35_9# Gnd 0.56fF
C1755 enable_0/2_input_AND_6/w_n12_9# Gnd 0.72fF
C1756 OUTPUT_ALU_ANDBLOCK_B1 Gnd 0.95fF
C1757 enable_0/2_input_AND_5/OUT Gnd 0.38fF
C1758 enable_0/2_input_AND_5/w_35_9# Gnd 0.56fF
C1759 enable_0/2_input_AND_5/w_n12_9# Gnd 0.72fF
C1760 OUTPUT_ALU_ANDBLOCK_B0 Gnd 0.90fF
C1761 enable_0/2_input_AND_4/OUT Gnd 0.38fF
C1762 enable_0/2_input_AND_4/w_35_9# Gnd 0.56fF
C1763 enable_0/2_input_AND_4/w_n12_9# Gnd 0.72fF
C1764 enable_0/2_input_AND_3/OUT Gnd 0.38fF
C1765 enable_0/2_input_AND_3/w_35_9# Gnd 0.56fF
C1766 enable_0/2_input_AND_3/w_n12_9# Gnd 0.72fF
C1767 enable_0/2_input_AND_2/OUT Gnd 0.38fF
C1768 enable_0/2_input_AND_2/w_35_9# Gnd 0.56fF
C1769 enable_0/2_input_AND_2/w_n12_9# Gnd 0.72fF
C1770 enable_0/2_input_AND_1/OUT Gnd 0.38fF
C1771 enable_0/2_input_AND_1/w_35_9# Gnd 0.56fF
C1772 enable_0/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1773 enable_0/2_input_AND_0/OUT Gnd 0.38fF
C1774 S0_S1_DECODER Gnd 4.66fF
C1775 enable_0/2_input_AND_0/w_35_9# Gnd 0.56fF
C1776 enable_0/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1777 OUTPUT_ALU_ANDBLOCK_B3 Gnd 1.09fF
C1778 enable_0/2_input_AND_7/OUT Gnd 0.38fF
C1779 enable_0/2_input_AND_7/w_35_9# Gnd 0.56fF
C1780 enable_0/2_input_AND_7/w_n12_9# Gnd 0.72fF
C1781 adder_subtractor_0/q1d_2_INPUT_XOR_4/ABAR Gnd 0.10fF
C1782 adder_subtractor_0/q1d_2_INPUT_XOR_4/BBAR Gnd 0.04fF
C1783 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_53_n17# Gnd 0.45fF
C1784 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_12_2# Gnd 0.04fF
C1785 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_n34_1# Gnd 0.08fF
C1786 adder_subtractor_0/q1d_2_INPUT_XOR_4/w_52_34# Gnd 0.45fF
C1787 adder_subtractor_0/q1d_2_INPUT_XOR_3/ABAR Gnd 0.10fF
C1788 adder_subtractor_0/q1d_2_INPUT_XOR_3/BBAR Gnd 0.04fF
C1789 OUTPUT_ALU_ADDER_B3 Gnd 0.95fF
C1790 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_53_n17# Gnd 0.45fF
C1791 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_12_2# Gnd 0.04fF
C1792 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_n34_1# Gnd 0.08fF
C1793 adder_subtractor_0/q1d_2_INPUT_XOR_3/w_52_34# Gnd 0.45fF
C1794 adder_subtractor_0/q1d_2_INPUT_XOR_2/ABAR Gnd 0.10fF
C1795 adder_subtractor_0/q1d_2_INPUT_XOR_2/BBAR Gnd 0.04fF
C1796 OUTPUT_ALU_ADDER_B2 Gnd 1.05fF
C1797 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_53_n17# Gnd 0.45fF
C1798 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_12_2# Gnd 0.04fF
C1799 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_n34_1# Gnd 0.08fF
C1800 adder_subtractor_0/q1d_2_INPUT_XOR_2/w_52_34# Gnd 0.45fF
C1801 adder_subtractor_0/q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C1802 adder_subtractor_0/q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C1803 OUTPUT_ALU_ADDER_B1 Gnd 1.08fF
C1804 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_53_n17# Gnd 0.45fF
C1805 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_12_2# Gnd 0.04fF
C1806 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_n34_1# Gnd 0.08fF
C1807 adder_subtractor_0/q1d_2_INPUT_XOR_1/w_52_34# Gnd 0.45fF
C1808 adder_subtractor_0/full_adder_3/2_input_AND_1/OUT Gnd 0.38fF
C1809 adder_subtractor_0/full_adder_3/AXORB Gnd 3.61fF
C1810 ADDER_SUB_C3 Gnd 2.57fF
C1811 adder_subtractor_0/full_adder_3/2_input_AND_1/w_35_9# Gnd 0.56fF
C1812 adder_subtractor_0/full_adder_3/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1813 adder_subtractor_0/full_adder_3/2_input_AND_0/OUT Gnd 0.38fF
C1814 OUTPUT_ALU_ADDER_A3 Gnd 2.38fF
C1815 adder_subtractor_0/full_adder_3/2_input_AND_0/w_35_9# Gnd 0.56fF
C1816 adder_subtractor_0/full_adder_3/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1817 ADDER_SUB_C4 Gnd 3.21fF
C1818 adder_subtractor_0/full_adder_3/2_input_OR_0/OUT Gnd 0.41fF
C1819 adder_subtractor_0/full_adder_3/2_input_OR_0/B Gnd 0.52fF
C1820 adder_subtractor_0/full_adder_3/2_input_OR_0/A Gnd 0.78fF
C1821 adder_subtractor_0/full_adder_3/2_input_OR_0/w_30_15# Gnd 0.60fF
C1822 adder_subtractor_0/full_adder_3/2_input_OR_0/w_n23_15# Gnd 0.73fF
C1823 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C1824 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C1825 ADDER_SUB_S3 Gnd 0.39fF
C1826 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_53_n17# Gnd 0.45fF
C1827 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_12_2# Gnd 0.04fF
C1828 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_n34_1# Gnd 0.08fF
C1829 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_1/w_52_34# Gnd 0.45fF
C1830 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1831 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1832 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1833 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1834 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1835 adder_subtractor_0/full_adder_3/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1836 adder_subtractor_0/full_adder_2/2_input_AND_1/OUT Gnd 0.38fF
C1837 adder_subtractor_0/full_adder_2/AXORB Gnd 3.61fF
C1838 ADDER_SUB_C2 Gnd 2.38fF
C1839 adder_subtractor_0/full_adder_2/2_input_AND_1/w_35_9# Gnd 0.56fF
C1840 adder_subtractor_0/full_adder_2/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1841 adder_subtractor_0/full_adder_2/2_input_AND_0/OUT Gnd 0.38fF
C1842 adder_subtractor_0/B2_XOR Gnd 4.17fF
C1843 OUTPUT_ALU_ADDER_A2 Gnd 2.32fF
C1844 adder_subtractor_0/full_adder_2/2_input_AND_0/w_35_9# Gnd 0.56fF
C1845 adder_subtractor_0/full_adder_2/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1846 adder_subtractor_0/full_adder_2/2_input_OR_0/OUT Gnd 0.41fF
C1847 adder_subtractor_0/full_adder_2/2_input_OR_0/B Gnd 0.52fF
C1848 adder_subtractor_0/full_adder_2/2_input_OR_0/A Gnd 0.78fF
C1849 adder_subtractor_0/full_adder_2/2_input_OR_0/w_30_15# Gnd 0.60fF
C1850 adder_subtractor_0/full_adder_2/2_input_OR_0/w_n23_15# Gnd 0.73fF
C1851 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C1852 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C1853 ADDER_SUB_S2 Gnd 0.31fF
C1854 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_53_n17# Gnd 0.45fF
C1855 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_12_2# Gnd 0.04fF
C1856 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_n34_1# Gnd 0.08fF
C1857 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_1/w_52_34# Gnd 0.45fF
C1858 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1859 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1860 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1861 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1862 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1863 adder_subtractor_0/full_adder_2/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1864 adder_subtractor_0/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1865 adder_subtractor_0/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1866 OUTPUT_ALU_ADDER_B0 Gnd 1.17fF
C1867 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1868 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1869 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1870 adder_subtractor_0/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1871 adder_subtractor_0/full_adder_1/2_input_AND_1/OUT Gnd 0.38fF
C1872 adder_subtractor_0/full_adder_1/AXORB Gnd 3.61fF
C1873 adder_subtractor_0/full_adder_1/2_input_AND_1/w_35_9# Gnd 0.56fF
C1874 adder_subtractor_0/full_adder_1/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1875 adder_subtractor_0/full_adder_1/2_input_AND_0/OUT Gnd 0.38fF
C1876 adder_subtractor_0/B1_XOR Gnd 3.96fF
C1877 OUTPUT_ALU_ADDER_A1 Gnd 2.32fF
C1878 adder_subtractor_0/full_adder_1/2_input_AND_0/w_35_9# Gnd 0.56fF
C1879 adder_subtractor_0/full_adder_1/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1880 adder_subtractor_0/full_adder_1/2_input_OR_0/OUT Gnd 0.41fF
C1881 adder_subtractor_0/full_adder_1/2_input_OR_0/B Gnd 0.52fF
C1882 adder_subtractor_0/full_adder_1/2_input_OR_0/A Gnd 0.78fF
C1883 adder_subtractor_0/full_adder_1/2_input_OR_0/w_30_15# Gnd 0.60fF
C1884 adder_subtractor_0/full_adder_1/2_input_OR_0/w_n23_15# Gnd 0.73fF
C1885 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C1886 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C1887 ADDER_SUB_S1 Gnd 0.33fF
C1888 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_53_n17# Gnd 0.45fF
C1889 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_12_2# Gnd 0.04fF
C1890 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_n34_1# Gnd 0.08fF
C1891 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_1/w_52_34# Gnd 0.45fF
C1892 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1893 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1894 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1895 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1896 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1897 adder_subtractor_0/full_adder_1/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1898 VDD Gnd 310.39fF
C1899 adder_subtractor_0/full_adder_0/2_input_AND_1/OUT Gnd 0.38fF
C1900 adder_subtractor_0/full_adder_0/AXORB Gnd 3.61fF
C1901 ADD_SUB_M Gnd 58.56fF
C1902 adder_subtractor_0/full_adder_0/2_input_AND_1/w_35_9# Gnd 0.56fF
C1903 adder_subtractor_0/full_adder_0/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1904 adder_subtractor_0/full_adder_0/2_input_AND_0/OUT Gnd 0.38fF
C1905 OUTPUT_ALU_ADDER_A0 Gnd 4.19fF
C1906 adder_subtractor_0/B0_XOR Gnd 2.78fF
C1907 adder_subtractor_0/full_adder_0/2_input_AND_0/w_35_9# Gnd 0.56fF
C1908 adder_subtractor_0/full_adder_0/2_input_AND_0/w_n12_9# Gnd 0.72fF
C1909 GND Gnd 410.31fF
C1910 adder_subtractor_0/full_adder_0/2_input_OR_0/OUT Gnd 0.41fF
C1911 adder_subtractor_0/full_adder_0/2_input_OR_0/B Gnd 0.52fF
C1912 adder_subtractor_0/full_adder_0/2_input_OR_0/A Gnd 0.78fF
C1913 adder_subtractor_0/full_adder_0/2_input_OR_0/w_30_15# Gnd 0.60fF
C1914 adder_subtractor_0/full_adder_0/2_input_OR_0/w_n23_15# Gnd 0.73fF
C1915 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/ABAR Gnd 0.10fF
C1916 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/BBAR Gnd 0.04fF
C1917 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_53_n17# Gnd 0.45fF
C1918 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_12_2# Gnd 0.04fF
C1919 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_n34_1# Gnd 0.08fF
C1920 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_1/w_52_34# Gnd 0.45fF
C1921 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C1922 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C1923 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C1924 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C1925 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C1926 adder_subtractor_0/full_adder_0/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C1927 AND_OUTPUT_A3B3 Gnd 0.11fF
C1928 and_block_0/2_input_AND_3/OUT Gnd 0.38fF
C1929 OUTPUT_ALU_ANDBLOCK_A3 Gnd 0.82fF
C1930 and_block_0/2_input_AND_3/w_35_9# Gnd 0.56fF
C1931 and_block_0/2_input_AND_3/w_n12_9# Gnd 0.72fF
C1932 AND_OUTPUT_A2B2 Gnd 0.16fF
C1933 and_block_0/2_input_AND_2/OUT Gnd 0.38fF
C1934 OUTPUT_ALU_ANDBLOCK_A2 Gnd 0.90fF
C1935 and_block_0/2_input_AND_2/w_35_9# Gnd 0.56fF
C1936 and_block_0/2_input_AND_2/w_n12_9# Gnd 0.72fF
C1937 AND_OUTPUT_A1B1 Gnd 0.16fF
C1938 and_block_0/2_input_AND_1/OUT Gnd 0.38fF
C1939 OUTPUT_ALU_ANDBLOCK_A1 Gnd 0.72fF
C1940 and_block_0/2_input_AND_1/w_35_9# Gnd 0.56fF
C1941 and_block_0/2_input_AND_1/w_n12_9# Gnd 0.72fF
C1942 AND_OUTPUT_A0B0 Gnd 0.16fF
C1943 and_block_0/2_input_AND_0/OUT Gnd 0.38fF
C1944 OUTPUT_ALU_ANDBLOCK_A0 Gnd 0.82fF
C1945 and_block_0/2_input_AND_0/w_35_9# Gnd 0.56fF
C1946 and_block_0/2_input_AND_0/w_n12_9# Gnd 0.72fF
.tran 1n 800n
*target text

.control
run
set color0 = rgb:f/f/e
set color1 = white
* plot v(S0_DECODER) v(S1_DECODER)+2
* plot v(S0BAR_S1BAR_DECODER) v(S0_S1BAR_DECODER)+2 v(S0BAR_S1_DECODER)+4 v(S0_S1_DECODER)+6
plot v(INPUT_ALU_A0) v(INPUT_ALU_A1)+2 v(INPUT_ALU_A2)+4 v(INPUT_ALU_A3)+6
plot v(INPUT_ALU_B0) v(INPUT_ALU_B1)+2 v(INPUT_ALU_B2)+4 v(INPUT_ALU_B3)+6
* plot v(OUTPUT_ALU_ANDBLOCK_A0) v(OUTPUT_ALU_ANDBLOCK_A1)+2 v(OUTPUT_ALU_ANDBLOCK_A2)+4 v(OUTPUT_ALU_ANDBLOCK_A3)+6
* plot v(OUTPUT_ALU_ANDBLOCK_B0) v(OUTPUT_ALU_ANDBLOCK_B1)+2 v(OUTPUT_ALU_ANDBLOCK_B2)+4 v(OUTPUT_ALU_ANDBLOCK_B3)+6
* plot v(OUTPUT_ALU_COMPARATOR_A0) v(OUTPUT_ALU_COMPARATOR_A1)+2 v(OUTPUT_ALU_COMPARATOR_A2)+4 v(OUTPUT_ALU_COMPARATOR_A3)+6
* plot v(OUTPUT_ALU_COMPARATOR_B0) v(OUTPUT_ALU_COMPARATOR_B1)+2 v(OUTPUT_ALU_COMPARATOR_B2)+4 v(OUTPUT_ALU_COMPARATOR_B3)+6
* plot v(OUTPUT_ALU_ADDER_A0) v(OUTPUT_ALU_ADDER_A1)+2 v(OUTPUT_ALU_ADDER_A2)+4 v(OUTPUT_ALU_ADDER_A3)+6
* plot v(OUTPUT_ALU_ADDER_B0) v(OUTPUT_ALU_ADDER_B1)+2 v(OUTPUT_ALU_ADDER_B2)+4 v(OUTPUT_ALU_ADDER_B3)+6
plot v(AND_OUTPUT_A0B0) v(AND_OUTPUT_A1B1)+2 v(AND_OUTPUT_A2B2)+4 v(AND_OUTPUT_A3B3)+6 
* plot v(COMPARATOR_A_EQUAL_B_FINAL) v(COMPARATOR_OUT_A_LESSTHAN_B)+2 v(COMPARATOR_OUT_A_GREATERTHAN_B)+4
* plot v(ADDER_SUB_S0) v(ADDER_SUB_S1)+2 v(ADDER_SUB_S2)+4 v(ADDER_SUB_S3)+6 v(ADDER_SUB_CFINAL)+8 
* plot v(ADD_SUB_M)
* plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6 
* plot v(B0) v(B1)+2 v(B2)+4 v(B3)+6
* plot v(node_c1) v(node_c2)+2 v(node_c3)+4 v(node_c4)+6 v(node_c_final)+8
* plot v(B0_XOR) v(B1_XOR)+2 v(B2_XOR)+4 v(B3_XOR)+6 
* plot v(SUM_0) v(SUM_1)+2 v(SUM_2)+4 v(SUM_3)+6 v(CARRY_FINAL)+8 
* plot v(CARRY_1) v(CARRY_2)+2 v(CARRY_3)+4 v(CARRY_4)+6 
* hardcopy image.ps v(S0) v(S1)+2 v(S2)+4 v(S3)+6 v(node_c_final)+8
quit
.end
.endc