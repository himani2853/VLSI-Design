magic
tech scmos
timestamp 1700257825
<< polycontact >>
rect -882 102 -860 112
rect -602 107 -584 118
rect -306 112 -288 123
rect 8 113 24 127
rect -1952 27 -1926 43
rect -1811 14 -1803 24
rect -1580 -1 -1565 14
rect -473 0 -460 6
rect -177 5 -164 10
rect 135 4 151 11
rect -753 -6 -741 0
rect -38 -76 -21 -63
rect 332 -75 342 -65
rect -1235 -98 -1217 -83
rect 103 -88 116 -77
rect -1091 -108 -1081 -97
rect -616 -99 -600 -89
rect -482 -107 -473 -97
rect -859 -175 -840 -163
rect -250 -171 -233 -160
rect -1780 -493 -1767 -484
rect -1658 -603 -1647 -595
<< metal1 >>
rect -895 136 372 166
rect -882 112 -860 136
rect -601 118 -585 136
rect -306 123 -290 136
rect 8 127 24 136
rect -1952 80 -1493 84
rect -690 84 -689 95
rect -1386 80 -1374 81
rect -1952 76 -1374 80
rect -1952 43 -1928 76
rect -1503 67 -1374 76
rect -1503 66 -1435 67
rect -1386 42 -1374 67
rect -750 52 -722 57
rect -1386 24 -1007 42
rect -1803 14 -1772 24
rect -1565 13 -1413 14
rect -1565 -1 -1411 13
rect -1566 -25 -1537 -20
rect -1446 -220 -1411 -1
rect -1237 -13 -1067 0
rect -1236 -83 -1217 -13
rect -1080 -24 -1067 -13
rect -1011 -9 -1007 24
rect -1011 -14 -915 -9
rect -753 -14 -741 -6
rect -920 -24 -915 -14
rect -728 -24 -722 52
rect -1080 -33 -938 -24
rect -920 -29 -722 -24
rect -950 -38 -938 -33
rect -950 -47 -857 -38
rect -1236 -97 -1235 -83
rect -714 -85 -689 84
rect -468 58 -408 63
rect -176 61 -141 66
rect -473 -13 -460 0
rect -416 -24 -408 58
rect -177 -2 -164 5
rect -541 -27 -408 -24
rect -549 -31 -408 -27
rect -150 -37 -141 61
rect -1081 -108 -1073 -97
rect -690 -99 -689 -85
rect -616 -49 -141 -37
rect -616 -89 -602 -49
rect -130 -62 -107 93
rect 330 85 372 136
rect 139 63 219 67
rect 135 -3 151 4
rect 205 -20 219 63
rect 142 -31 219 -20
rect 330 62 611 85
rect -108 -71 -107 -62
rect -38 -63 -22 -32
rect 330 -65 372 62
rect 330 -73 332 -65
rect 342 -73 372 -65
rect 116 -87 128 -78
rect 116 -88 140 -87
rect -616 -100 -602 -99
rect -473 -107 -443 -97
rect 348 -127 392 -122
rect -848 -148 -823 -143
rect -240 -150 -216 -145
rect -840 -175 -720 -164
rect -233 -171 -138 -160
rect -1446 -244 -1410 -220
rect -1657 -301 -1646 -300
rect -1667 -305 -1646 -301
rect -1657 -384 -1646 -305
rect -1445 -317 -1410 -244
rect -1780 -397 -1646 -384
rect -1446 -363 -1410 -317
rect -1780 -484 -1767 -397
rect -1446 -449 -1411 -363
rect -949 -428 -928 -424
rect -1448 -466 -1411 -449
rect -933 -466 -928 -428
rect -1448 -471 -928 -466
rect -1448 -472 -1078 -471
rect -743 -476 -720 -175
rect -337 -430 -311 -426
rect -321 -476 -311 -430
rect -152 -454 -138 -171
rect 265 -403 276 -402
rect 247 -407 276 -403
rect 265 -454 276 -407
rect -152 -466 276 -454
rect -743 -483 -311 -476
rect 553 -512 611 62
rect -1655 -543 -1609 -536
rect 553 -569 612 -512
rect -1658 -607 -1648 -603
rect -1658 -608 -1216 -607
rect 556 -608 612 -569
rect -1658 -634 612 -608
rect -1290 -635 612 -634
<< m2contact >>
rect -816 88 -809 96
rect -864 82 -857 87
rect -714 84 -690 98
rect -582 88 -575 96
rect -533 90 -524 97
rect -292 90 -283 97
rect -241 94 -235 100
rect -130 93 -106 104
rect 26 94 32 100
rect -864 21 -858 26
rect -817 16 -812 21
rect -857 -47 -832 -36
rect -581 27 -575 32
rect -533 22 -528 27
rect -550 -27 -541 -15
rect -288 32 -283 38
rect -241 25 -236 31
rect -714 -99 -690 -85
rect 27 32 32 38
rect 74 26 81 32
rect 128 -31 142 -20
rect -132 -73 -108 -62
rect 128 -87 141 -75
rect -1767 -515 -1761 -507
rect -1720 -579 -1712 -573
<< metal2 >>
rect -1326 141 -1292 143
rect -2047 112 -1292 141
rect -2044 20 -2020 112
rect -1326 105 -1292 112
rect -1326 87 -917 105
rect -809 88 -714 96
rect -1326 83 -864 87
rect -1325 82 -864 83
rect -690 88 -582 96
rect -524 90 -292 97
rect -235 94 -130 100
rect -106 94 26 100
rect -1325 81 -955 82
rect -1323 -98 -1300 81
rect -299 32 -288 38
rect 15 32 27 37
rect -948 26 -915 30
rect -590 27 -581 32
rect -357 27 -340 28
rect -299 27 -293 32
rect 15 31 21 32
rect -948 21 -864 26
rect -948 17 -915 21
rect -945 -64 -920 17
rect -590 20 -585 27
rect -528 22 -293 27
rect -236 25 21 31
rect 81 26 433 32
rect -812 16 -585 20
rect -651 -27 -550 -15
rect -651 -37 -643 -27
rect -832 -47 -643 -37
rect -357 -59 -340 22
rect -947 -72 -759 -64
rect -357 -71 -152 -59
rect -783 -92 -759 -72
rect -174 -94 -152 -71
rect 128 -75 141 -31
rect 412 -73 433 26
rect -1921 -506 -1891 -265
rect -1504 -351 -1484 -312
rect -1505 -391 -1482 -351
rect -1507 -498 -1482 -391
rect -1921 -514 -1767 -506
rect -1507 -507 -1484 -498
rect -787 -507 -762 -429
rect -1507 -524 -762 -507
rect -1509 -536 -762 -524
rect -1509 -538 -764 -536
rect -1720 -585 -1713 -579
rect -1509 -585 -1470 -538
rect -1720 -594 -1469 -585
use q1d_2_INPUT_XOR  q1d_2_INPUT_XOR_0
timestamp 1699251415
transform 1 0 56 0 1 62
box -56 -62 103 58
use q1d_2_INPUT_XOR  q1d_2_INPUT_XOR_1
timestamp 1699251415
transform 1 0 -259 0 1 61
box -56 -62 103 58
use q1d_2_INPUT_XOR  q1d_2_INPUT_XOR_2
timestamp 1699251415
transform 1 0 -551 0 1 57
box -56 -62 103 58
use q1d_2_INPUT_XOR  q1d_2_INPUT_XOR_3
timestamp 1699251415
transform 1 0 -834 0 1 51
box -56 -62 103 58
use full_adder  full_adder_0
timestamp 1699686506
transform 1 0 -11 0 1 -218
box -119 -217 443 160
use full_adder  full_adder_1
timestamp 1699686506
transform 1 0 -596 0 1 -241
box -119 -217 443 160
use full_adder  full_adder_2
timestamp 1699686506
transform 1 0 -1205 0 1 -239
box -119 -217 443 160
use full_adder  full_adder_3
timestamp 1699686506
transform 1 0 -1925 0 1 -116
box -119 -217 443 160
use q1d_2_INPUT_XOR  q1d_2_INPUT_XOR_4
timestamp 1699251415
transform 1 0 -1738 0 1 -544
box -56 -62 103 58
<< labels >>
rlabel metal1 -63 149 -58 152 1 M
rlabel metal1 141 -2 142 -1 1 B0
rlabel metal1 164 64 165 65 7 B0_XOR
rlabel metal1 -170 0 -170 1 1 B1
rlabel metal1 -148 62 -147 63 1 B1_XOR
rlabel metal1 -467 -10 -466 -8 1 B2
rlabel metal1 -440 59 -438 61 1 B2_XOR
rlabel metal1 -748 -10 -746 -9 1 B3
rlabel metal1 -726 54 -724 55 1 B3_XOR
rlabel metal2 -940 94 -936 97 1 VDD
rlabel metal2 -935 23 -933 24 1 GND
rlabel metal1 -31 -47 -30 -40 1 A0
rlabel metal1 378 -125 381 -124 1 SUM_0
rlabel metal1 263 -406 264 -405 1 CARRY_1
rlabel metal1 -455 -105 -449 -103 1 A1
rlabel metal1 -221 -148 -220 -147 1 SUM_1
rlabel metal1 -328 -429 -326 -427 1 CARRY_2
rlabel metal1 -1078 -102 -1077 -101 1 A2
rlabel metal1 -828 -146 -827 -145 1 SUM_2
rlabel metal1 -936 -426 -933 -425 1 CARRY_3
rlabel metal1 -1785 19 -1783 22 1 A3
rlabel metal1 -1544 -24 -1543 -22 1 SUM_3
rlabel metal1 -1656 -303 -1654 -302 1 CARRY_4
rlabel metal1 -1619 -540 -1614 -538 1 CARRY_FINAL
<< end >>
