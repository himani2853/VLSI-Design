.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include OR.sub
.include XNOR.sub
.include XOR.sub
.include 4_input_AND.sub
.include 4_input_OR.sub
.include 3_input_AND.sub
.include 5_input_AND.sub
.include comparator.sub


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 node_a0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)
* V_in_c node_m gnd PULSE(0 1.8 0ns 100ps 100ps 400ns 800ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)

* V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 100ns 160ns)
* V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 200ns 240ns)
* V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 400ns 520ns)
* V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 600ns 800ns)

X1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_equal_final node_ALB_final node_AGB_final node_x gnd comparator


.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a0) v(node_a1)+2 v(node_a2)+4 v(node_a3)+6 v(node_b0)+8 v(node_b1)+10 v(node_b2)+12 v(node_b3)+14
plot v(node_ALB_final) v(node_equal_final)+2 v(node_AGB_final)+4
* hardcopy image.ps v(node_a0) v(node_a1)+2 v(node_a2)+4 v(node_a3)+6
.end
.endc