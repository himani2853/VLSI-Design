magic
tech scmos
timestamp 1701471188
<< metal1 >>
rect 4106 1418 4158 1423
rect 3526 1412 4158 1418
rect 1709 1397 4158 1412
rect -79 1395 536 1396
rect 885 1395 4158 1397
rect -79 1381 4158 1395
rect -79 1358 13 1381
rect 30 1378 4158 1381
rect 30 1362 1141 1378
rect 30 1358 912 1362
rect -513 1310 -285 1311
rect -513 1308 -37 1310
rect -513 1307 320 1308
rect -513 1302 438 1307
rect -513 1301 320 1302
rect -513 1300 -37 1301
rect -513 1123 -496 1300
rect 433 1276 437 1302
rect 486 1281 498 1358
rect 525 1356 912 1358
rect 434 1199 437 1203
rect 430 1195 437 1199
rect 434 1180 438 1195
rect -513 1071 -494 1123
rect 433 1098 435 1102
rect 442 1101 445 1106
rect 432 1095 439 1098
rect 435 1077 439 1095
rect -512 724 -494 1071
rect 442 1000 446 1004
rect 432 996 439 998
rect 427 994 439 996
rect 435 979 439 994
rect 432 903 433 908
rect 429 900 439 903
rect 436 899 439 900
rect 436 886 440 899
rect 428 803 432 805
rect 428 800 441 803
rect 437 780 441 800
rect -514 447 -494 724
rect 430 696 442 699
rect 438 675 442 696
rect 351 602 365 612
rect 445 602 449 605
rect 351 583 359 602
rect 435 592 439 599
rect 445 597 453 602
rect 435 591 445 592
rect 435 589 454 591
rect 442 588 454 589
rect 315 582 359 583
rect 98 573 359 582
rect 449 574 454 588
rect 99 487 103 573
rect 351 572 359 573
rect 441 570 454 574
rect 381 520 392 542
rect 99 483 114 487
rect 99 469 103 483
rect 380 474 392 520
rect 448 493 452 495
rect 380 464 391 474
rect -514 441 -503 447
rect 186 441 187 445
rect 205 441 451 445
rect -514 171 -496 441
rect 447 407 451 441
rect 572 431 600 1356
rect 648 1323 674 1356
rect 919 1361 1141 1362
rect 1156 1361 4158 1378
rect 919 1359 4158 1361
rect 919 1356 930 1359
rect 1709 1357 4158 1359
rect 3689 1355 4158 1357
rect 648 1158 672 1323
rect 648 1117 673 1158
rect 649 544 673 1117
rect 857 1109 867 1113
rect 863 1094 867 1109
rect 879 1014 890 1018
rect 862 1001 866 1012
rect 879 925 890 929
rect 862 908 866 918
rect 862 830 863 834
rect 880 832 891 836
rect 862 817 866 830
rect 869 816 873 819
rect 876 738 896 742
rect 856 628 1144 629
rect 856 627 1916 628
rect 856 625 2331 627
rect 856 624 2304 625
rect 855 613 2304 624
rect 649 514 674 544
rect 500 414 600 431
rect 501 399 513 414
rect 90 361 93 367
rect 237 364 351 365
rect 178 360 351 364
rect 362 360 376 365
rect 178 359 376 360
rect 650 348 674 514
rect 855 470 870 613
rect 1901 612 2304 613
rect 902 589 916 590
rect 901 588 1088 589
rect 901 587 1278 588
rect 1473 587 1989 590
rect 901 579 1989 587
rect 902 518 916 579
rect 795 465 870 470
rect -400 329 -50 333
rect 572 330 630 335
rect 442 327 451 329
rect 442 326 452 327
rect 448 312 452 326
rect 649 308 674 348
rect 794 458 870 465
rect 165 261 176 265
rect 583 233 631 239
rect 443 226 453 229
rect 23 219 38 223
rect 449 209 453 226
rect -516 -225 -496 171
rect 649 163 673 308
rect 565 130 635 137
rect 446 125 453 128
rect 449 112 453 125
rect 648 112 673 163
rect 32 -70 35 61
rect 451 33 453 37
rect 566 33 630 38
rect 450 28 453 33
rect 450 18 454 28
rect 104 -9 108 18
rect 104 -12 116 -9
rect 104 -15 108 -12
rect 52 -21 108 -15
rect 52 -24 57 -21
rect 52 -63 57 -29
rect 648 -44 672 112
rect 794 44 806 458
rect 855 457 870 458
rect 903 398 916 518
rect 1039 540 1050 541
rect 1039 530 1040 540
rect 3104 532 3110 660
rect 4106 577 4158 1355
rect 3208 563 4158 577
rect 3207 535 3222 539
rect 1039 478 1050 530
rect 3104 528 3138 532
rect 3052 521 3140 525
rect 3203 509 3427 517
rect 3398 490 3427 509
rect 1038 457 1050 478
rect 1038 403 1049 457
rect 2405 432 2413 433
rect 1989 431 1996 432
rect 903 366 917 398
rect 1038 394 1050 403
rect 1989 396 1996 421
rect 2405 406 2413 425
rect 2873 402 2886 407
rect 904 140 917 366
rect 1039 241 1050 394
rect 2533 310 2586 314
rect 2533 309 2538 310
rect 1304 301 1329 306
rect 1304 291 1310 301
rect 1738 297 1761 304
rect 2144 301 2186 305
rect 2537 305 2538 309
rect 2144 298 2149 301
rect 1309 283 1310 291
rect 2144 290 2149 291
rect 1154 213 1174 232
rect 916 130 917 140
rect 2488 162 2532 172
rect 2488 161 2540 162
rect 2488 80 2495 161
rect 2487 64 2495 80
rect 2487 53 2494 64
rect 2486 23 2494 53
rect 2486 4 2493 23
rect 2486 -4 2525 4
rect 1128 -18 1141 -17
rect 1128 -29 1269 -18
rect 52 -67 89 -63
rect 446 -64 449 -59
rect 547 -61 629 -57
rect 445 -68 455 -64
rect 32 -74 101 -70
rect 161 -74 232 -68
rect 221 -135 231 -74
rect 451 -87 455 -68
rect 648 -73 673 -44
rect -516 -407 -498 -225
rect 80 -304 107 -148
rect -516 -416 -25 -407
rect -495 -417 -25 -416
rect 81 -411 107 -304
rect -495 -418 -14 -417
rect 220 -448 231 -135
rect 581 -165 630 -160
rect 458 -190 461 -175
rect 452 -193 461 -190
rect 561 -271 635 -266
rect 644 -271 645 -266
rect 451 -276 468 -273
rect 464 -294 468 -276
rect 455 -298 468 -294
rect 341 -378 343 -355
rect 371 -378 405 -355
rect 341 -379 405 -378
rect 462 -382 633 -378
rect 281 -402 463 -399
rect 220 -460 389 -448
rect 459 -463 463 -402
rect 649 -456 673 -73
rect 1128 -117 1141 -29
rect 1294 -29 1297 -18
rect 1070 -118 1141 -117
rect 1079 -128 1141 -118
rect 2509 -209 2523 -4
rect 2872 -102 2887 -76
rect 1286 -265 1298 -262
rect 1382 -254 1573 -253
rect 1382 -262 1996 -254
rect 1541 -263 1996 -262
rect 1029 -271 1298 -265
rect 1029 -272 1296 -271
rect 1211 -332 1327 -321
rect 1314 -364 1327 -332
rect 2508 -362 2524 -209
rect 2465 -363 2524 -362
rect 2388 -364 2524 -363
rect 1314 -365 1682 -364
rect 2178 -365 2524 -364
rect 1314 -366 1766 -365
rect 1945 -366 2524 -365
rect 1314 -374 2524 -366
rect 1314 -378 2523 -374
rect 1314 -379 2432 -378
rect 1314 -380 2347 -379
rect 2465 -380 2523 -378
rect 1597 -381 2186 -380
rect 1753 -382 2017 -381
rect 512 -482 673 -456
rect -513 -538 139 -519
rect -513 -543 135 -538
rect 461 -542 463 -539
rect -513 -545 139 -543
rect 460 -545 463 -542
rect 460 -560 464 -545
rect 228 -643 366 -636
rect 229 -683 248 -643
rect 455 -644 465 -641
rect 461 -660 465 -644
rect -547 -714 248 -683
rect 456 -742 460 -740
rect 456 -745 465 -742
rect -515 -755 -11 -747
rect -515 -756 -94 -755
rect 461 -759 465 -745
rect 463 -835 465 -831
rect 462 -840 465 -835
rect 462 -853 466 -840
rect 598 -931 761 -927
rect 455 -938 474 -935
rect 471 -952 474 -938
rect 463 -956 474 -952
rect 698 -1031 705 -1030
rect 586 -1035 705 -1031
rect 465 -1042 474 -1038
rect 470 -1061 474 -1042
rect 464 -1065 474 -1061
rect 639 -1135 644 -1134
rect 572 -1140 644 -1135
rect 464 -1148 479 -1145
rect 475 -1165 479 -1148
rect 639 -1164 644 -1140
rect 467 -1168 479 -1165
rect 4 -1465 32 -1441
rect 66 -1465 81 -1441
rect 4 -1470 81 -1465
rect 406 -1441 418 -1231
rect 474 -1259 478 -1243
rect 637 -1253 645 -1164
rect 2144 -1165 2164 -1157
rect 637 -1260 646 -1253
rect 638 -1302 646 -1260
rect 638 -1349 647 -1302
rect 639 -1371 647 -1349
rect 2838 -1436 3240 -1433
rect 734 -1441 3240 -1436
rect 117 -1467 602 -1441
rect 631 -1467 3240 -1441
rect 117 -1469 3240 -1467
rect 117 -1470 3042 -1469
rect 734 -1472 3042 -1470
rect 734 -1473 1508 -1472
rect 2063 -1518 2081 -1472
rect 3399 -1433 3425 490
rect 3312 -1458 3573 -1433
rect 3724 -1458 4026 -1429
rect 3312 -1469 4026 -1458
rect 3399 -1470 3425 -1469
rect 3677 -1472 4026 -1469
rect 2064 -1551 2080 -1518
rect 665 -1567 970 -1566
rect 1046 -1567 1303 -1566
rect -28 -1568 340 -1567
rect 665 -1568 1829 -1567
rect 2287 -1568 2313 -1567
rect -28 -1569 2060 -1568
rect 2226 -1569 2313 -1568
rect -28 -1592 2313 -1569
rect -28 -1593 1177 -1592
rect 1232 -1593 2313 -1592
rect -28 -1594 970 -1593
rect 1803 -1594 2313 -1593
rect -28 -1595 688 -1594
rect 2013 -1595 2313 -1594
rect 4106 -1577 4158 563
rect 2727 -1580 4158 -1577
rect 2522 -1593 4158 -1580
rect 309 -1596 688 -1595
rect 2226 -1598 2313 -1595
rect 2064 -1659 2079 -1610
rect 2287 -1652 2313 -1598
rect 2130 -1659 2257 -1658
rect 2064 -1675 2257 -1659
rect 2064 -1676 2191 -1675
rect 2249 -1757 2257 -1675
rect 2287 -1682 2368 -1652
rect 3595 -1673 3662 -1660
rect 2249 -1765 2291 -1757
rect 2282 -1788 2291 -1765
rect 2573 -1828 2586 -1717
rect 2573 -1831 2770 -1828
rect 2478 -1832 2490 -1831
rect 2475 -1838 2490 -1832
rect 2853 -1834 2860 -1710
rect 3054 -1833 3068 -1819
rect 2977 -1834 3069 -1833
rect 1685 -1844 1708 -1839
rect 2853 -1840 3069 -1834
rect 2977 -1842 3069 -1840
rect 3179 -1851 3188 -1706
rect 3210 -1825 3215 -1711
rect 3366 -1825 3382 -1818
rect 3210 -1828 3382 -1825
rect 3179 -1857 3209 -1851
rect 3606 -1946 3692 -1941
rect 2400 -1966 2417 -1961
rect 3012 -1969 3022 -1964
rect 1582 -2131 1610 -2121
rect 3499 -2226 3523 -2220
rect 2300 -2249 2317 -2245
rect 2915 -2257 2940 -2251
rect 1620 -2362 1634 -2355
<< m2contact >>
rect 13 1353 30 1381
rect 428 1199 434 1204
rect 442 1198 447 1203
rect 427 1098 433 1103
rect 445 1100 450 1106
rect 427 996 432 1002
rect 446 1000 451 1005
rect 426 903 432 908
rect 444 902 449 907
rect 426 805 432 810
rect 443 806 449 812
rect 429 699 434 704
rect 444 702 451 710
rect 365 602 374 612
rect 430 594 435 599
rect 453 595 461 603
rect 448 484 455 493
rect 380 452 394 464
rect -503 441 -493 447
rect 187 441 205 446
rect 912 1353 919 1362
rect 1141 1361 1156 1378
rect 851 1108 857 1116
rect 870 1093 875 1098
rect 862 1012 868 1017
rect 869 1002 874 1008
rect 857 913 862 919
rect 869 907 874 913
rect 863 830 868 835
rect 869 819 874 824
rect 3098 660 3111 683
rect 99 359 104 364
rect 172 359 178 365
rect 351 360 362 370
rect 376 359 387 365
rect 2304 612 2334 625
rect 1989 579 1996 590
rect -436 327 -400 337
rect -50 327 -32 334
rect 442 329 447 334
rect 454 330 460 335
rect 563 330 572 336
rect 630 330 641 336
rect 440 229 447 234
rect 455 233 462 240
rect 572 233 583 239
rect 631 233 639 241
rect 445 128 450 133
rect 456 131 462 137
rect 554 130 565 137
rect 635 130 644 138
rect 97 108 102 113
rect 31 61 36 67
rect 446 33 451 38
rect 456 33 462 38
rect 557 33 566 39
rect 630 33 639 38
rect 51 -29 58 -24
rect 1040 530 1054 540
rect 3039 519 3052 525
rect 1141 479 1152 488
rect 1989 421 1996 431
rect 1566 396 1576 408
rect 2405 425 2413 432
rect 2886 400 2896 408
rect 1116 330 1127 337
rect 1729 297 1738 305
rect 2532 304 2537 309
rect 2143 291 2150 298
rect 1303 282 1309 291
rect 1039 232 1050 241
rect 2897 196 2923 225
rect 904 130 916 140
rect 2532 162 2541 176
rect 794 33 807 44
rect 439 -64 446 -59
rect 457 -61 463 -56
rect 540 -61 547 -56
rect 629 -61 634 -56
rect 79 -148 111 -126
rect -25 -417 -10 -405
rect 81 -434 107 -411
rect 458 -165 463 -160
rect 570 -165 581 -159
rect 630 -165 637 -159
rect 457 -175 462 -170
rect 459 -270 464 -265
rect 550 -271 561 -265
rect 446 -276 451 -271
rect 635 -272 644 -264
rect 343 -378 371 -353
rect 633 -382 643 -377
rect 272 -402 281 -397
rect 389 -460 402 -447
rect 1269 -30 1294 -16
rect 1070 -128 1079 -118
rect 1284 -262 1299 -251
rect 1356 -263 1382 -253
rect 1996 -263 2010 -254
rect 1019 -272 1029 -265
rect 1198 -334 1211 -319
rect -541 -545 -513 -519
rect 135 -543 140 -538
rect 456 -542 461 -537
rect 468 -541 476 -533
rect 467 -636 475 -629
rect 366 -643 373 -636
rect 455 -641 460 -636
rect -575 -714 -547 -679
rect 455 -740 460 -735
rect 468 -739 475 -734
rect -547 -759 -515 -742
rect -11 -756 0 -747
rect 458 -835 463 -830
rect 468 -837 473 -832
rect 469 -931 475 -926
rect 592 -931 598 -926
rect 450 -938 455 -933
rect 761 -934 772 -924
rect 470 -1035 475 -1030
rect 576 -1035 586 -1028
rect 705 -1037 735 -1030
rect 460 -1042 465 -1037
rect 471 -1140 477 -1135
rect 565 -1140 572 -1135
rect 459 -1148 464 -1143
rect 32 -1465 66 -1431
rect 81 -1470 117 -1433
rect 473 -1265 479 -1259
rect 639 -1403 651 -1371
rect 602 -1467 631 -1441
rect 3240 -1477 3312 -1423
rect 3573 -1458 3724 -1427
rect 2064 -1559 2081 -1551
rect -50 -1595 -28 -1562
rect 2506 -1595 2522 -1576
rect 2063 -1610 2080 -1600
rect 2573 -1717 2587 -1704
rect 2853 -1710 2861 -1698
rect 3179 -1706 3188 -1698
rect 1449 -1805 1460 -1794
rect 2282 -1803 2294 -1788
rect 2468 -1838 2475 -1832
rect 3210 -1711 3215 -1703
rect 2153 -1927 2164 -1914
rect 2777 -1927 2788 -1915
<< metal2 >>
rect 15 1158 27 1353
rect 405 1199 428 1204
rect 447 1198 874 1203
rect -659 1105 -622 1106
rect -659 1095 -387 1105
rect -659 1093 -356 1095
rect -659 1092 -622 1093
rect -789 992 -458 1007
rect -88 774 -73 832
rect -265 699 -259 712
rect -241 699 -239 712
rect -265 564 -239 699
rect -179 572 -153 741
rect -86 686 -73 774
rect -89 574 -70 686
rect 15 668 26 1158
rect 852 1116 857 1139
rect 410 1098 427 1102
rect 445 1094 827 1100
rect 820 1028 827 1094
rect 870 1098 874 1198
rect 912 1096 918 1353
rect 1142 1290 1156 1361
rect 858 1012 862 1017
rect 410 1002 432 1003
rect 410 996 427 1002
rect 874 1002 878 1023
rect 446 998 451 1000
rect 446 994 760 998
rect 560 993 760 994
rect 755 966 760 993
rect 755 965 807 966
rect 755 960 820 965
rect 814 939 819 960
rect 857 919 862 921
rect 869 913 877 919
rect 407 903 426 908
rect 449 902 749 906
rect 444 899 749 902
rect 745 873 749 899
rect 745 866 802 873
rect 797 847 802 866
rect 859 830 863 834
rect 874 820 878 840
rect 411 805 426 810
rect 449 806 574 811
rect 835 726 842 756
rect 411 699 429 704
rect 451 702 623 708
rect 835 697 3731 726
rect 1260 673 3098 683
rect 1107 672 3098 673
rect -493 441 -21 447
rect 15 380 25 668
rect 1115 662 3098 672
rect 1260 660 3098 662
rect 2334 624 2393 625
rect 2334 612 2396 624
rect 407 594 430 599
rect 461 595 690 599
rect 453 594 690 595
rect 1054 530 1577 540
rect 690 492 772 493
rect 455 484 772 492
rect 1141 488 1151 498
rect 1566 504 1577 530
rect 1989 527 1996 579
rect 615 462 626 463
rect 394 452 626 462
rect 165 441 187 446
rect 351 370 361 432
rect 615 416 626 452
rect 1989 431 1995 446
rect 2405 432 2413 439
rect 613 410 626 416
rect 104 359 172 364
rect 178 359 179 364
rect -573 327 -436 334
rect -400 327 -396 334
rect -32 329 -25 333
rect 394 329 442 333
rect 460 330 563 335
rect 613 298 625 410
rect 1566 408 1576 422
rect 3039 407 3052 519
rect 2896 400 3052 407
rect 3039 399 3052 400
rect 749 335 1116 336
rect 641 330 1116 335
rect 612 289 625 298
rect 1711 297 1729 304
rect 2537 304 2538 307
rect 1711 292 1719 297
rect -647 233 -52 246
rect 422 230 440 234
rect 462 233 572 239
rect 612 191 624 289
rect 1295 283 1303 290
rect 1309 283 1310 290
rect 2092 291 2093 297
rect 2107 291 2143 297
rect 2532 243 2538 304
rect 639 239 748 240
rect 639 238 926 239
rect 639 233 1039 238
rect 720 232 1039 233
rect 1050 232 1052 238
rect 2531 211 2538 243
rect 3242 225 3307 226
rect 2531 202 2539 211
rect -768 158 -54 175
rect 611 171 624 191
rect 2532 176 2539 202
rect 2923 196 3307 225
rect 420 128 445 132
rect 462 131 554 137
rect 51 108 97 112
rect 51 89 55 108
rect 32 84 55 89
rect 32 67 35 84
rect 423 33 446 37
rect 462 33 557 38
rect 244 10 256 12
rect 191 0 256 10
rect 8 -24 21 -23
rect 8 -25 51 -24
rect 7 -28 51 -25
rect -105 -72 -35 -54
rect -105 -73 -20 -72
rect 7 -79 19 -28
rect 8 -96 19 -79
rect 8 -116 20 -96
rect 9 -129 20 -116
rect 7 -135 20 -129
rect -231 -161 -120 -160
rect -231 -162 -112 -161
rect -231 -180 -29 -162
rect -244 -181 -112 -180
rect -325 -244 -24 -219
rect -346 -245 -24 -244
rect 7 -265 19 -135
rect 244 -127 256 0
rect 422 -64 439 -59
rect 463 -61 540 -57
rect 111 -148 256 -127
rect 244 -149 256 -148
rect 413 -170 416 -164
rect 463 -165 570 -161
rect 413 -173 457 -170
rect -52 -279 19 -265
rect 464 -270 550 -266
rect 420 -276 446 -273
rect -53 -281 19 -279
rect -53 -402 -40 -281
rect 33 -352 68 -350
rect 27 -353 205 -352
rect 27 -378 343 -353
rect 27 -379 369 -378
rect 27 -380 205 -379
rect -53 -498 -39 -402
rect -10 -416 1 -405
rect -10 -417 3 -416
rect 33 -476 68 -380
rect 174 -402 272 -399
rect 174 -410 181 -402
rect -53 -502 -37 -498
rect -575 -544 -541 -519
rect -52 -644 -37 -502
rect -50 -664 -37 -644
rect 29 -522 68 -476
rect 80 -411 107 -410
rect 80 -434 81 -411
rect -648 -712 -575 -684
rect -50 -740 -36 -664
rect -767 -757 -547 -748
rect -49 -1075 -36 -740
rect 0 -755 8 -747
rect 29 -917 63 -522
rect 80 -917 107 -434
rect 611 -438 622 171
rect 644 130 904 137
rect 699 38 794 40
rect 639 33 794 38
rect 807 33 808 40
rect 1294 -29 1305 -19
rect 1294 -30 1324 -29
rect 684 -57 1071 -55
rect 634 -61 1071 -57
rect 684 -62 1071 -61
rect 1071 -159 1078 -128
rect 739 -160 1079 -159
rect 637 -165 1079 -160
rect 1299 -262 1356 -253
rect 1382 -262 1383 -253
rect 2010 -256 2050 -255
rect 2010 -262 2024 -256
rect 2010 -263 2050 -262
rect 644 -272 1019 -266
rect 1195 -334 1198 -320
rect 1195 -376 1210 -334
rect 3242 -346 3307 196
rect 909 -378 1210 -376
rect 643 -382 1210 -378
rect 909 -383 1200 -382
rect 140 -543 146 -539
rect 431 -542 456 -539
rect 476 -540 580 -533
rect 611 -612 624 -438
rect 373 -643 377 -636
rect 475 -636 586 -632
rect 429 -641 455 -636
rect 434 -740 455 -736
rect 475 -739 558 -735
rect 427 -835 458 -831
rect 473 -837 565 -834
rect -50 -1104 -36 -1075
rect -50 -1281 -37 -1104
rect -50 -1317 -36 -1281
rect -49 -1498 -36 -1317
rect 29 -1431 63 -921
rect 29 -1452 32 -1431
rect 80 -1433 107 -921
rect 425 -935 429 -921
rect 475 -931 592 -928
rect 425 -938 450 -935
rect 613 -1017 624 -612
rect 475 -1035 576 -1031
rect 439 -1042 460 -1038
rect 477 -1140 565 -1136
rect 431 -1148 459 -1145
rect 474 -1259 478 -1258
rect 80 -1464 81 -1433
rect -50 -1562 -33 -1498
rect 474 -1617 478 -1265
rect 612 -1440 624 -1017
rect 638 -1403 639 -1374
rect 705 -1390 733 -1037
rect 761 -1046 772 -934
rect 761 -1065 771 -1046
rect 759 -1088 771 -1065
rect 758 -1291 771 -1088
rect 3240 -1177 3307 -346
rect 3239 -1239 3307 -1177
rect 758 -1330 769 -1291
rect 758 -1342 768 -1330
rect 3146 -1341 3158 -1340
rect 1368 -1342 3158 -1341
rect 758 -1352 3158 -1342
rect 758 -1353 1381 -1352
rect 3146 -1369 3158 -1352
rect 2352 -1382 2663 -1381
rect 2227 -1383 2663 -1382
rect 2100 -1384 2663 -1383
rect 1975 -1385 2663 -1384
rect 1925 -1386 2663 -1385
rect 1839 -1387 2663 -1386
rect 1711 -1388 2663 -1387
rect 1649 -1389 2663 -1388
rect 896 -1390 2663 -1389
rect 705 -1399 2663 -1390
rect 705 -1400 2415 -1399
rect 705 -1401 2270 -1400
rect 705 -1402 2161 -1401
rect 705 -1403 2020 -1402
rect 610 -1441 625 -1440
rect 638 -1493 646 -1403
rect 705 -1404 1989 -1403
rect 705 -1405 1460 -1404
rect 1581 -1405 1867 -1404
rect 705 -1406 733 -1405
rect 1581 -1406 1744 -1405
rect 1581 -1407 1676 -1406
rect 636 -1524 648 -1493
rect 2645 -1511 2663 -1399
rect 2853 -1509 2860 -1508
rect 2789 -1510 2861 -1509
rect 2720 -1511 2861 -1510
rect 2645 -1523 2861 -1511
rect 2645 -1524 2791 -1523
rect 635 -1530 649 -1524
rect 2645 -1526 2663 -1524
rect 2059 -1528 2339 -1527
rect 1993 -1529 2339 -1528
rect 993 -1530 1238 -1529
rect 1567 -1530 2339 -1529
rect 635 -1532 1396 -1530
rect 1414 -1531 2537 -1530
rect 1414 -1532 2587 -1531
rect 635 -1543 2587 -1532
rect 642 -1544 2587 -1543
rect 993 -1545 2587 -1544
rect 1151 -1546 1659 -1545
rect 1285 -1548 1530 -1546
rect 1673 -1547 1918 -1545
rect 1993 -1546 2587 -1545
rect 1993 -1547 2158 -1546
rect 2271 -1549 2587 -1546
rect 1448 -1652 1459 -1564
rect 2064 -1600 2079 -1559
rect 2153 -1655 2166 -1561
rect 2291 -1593 2506 -1580
rect 1449 -1794 1459 -1726
rect 2291 -1731 2301 -1593
rect 2573 -1606 2587 -1549
rect 2573 -1704 2586 -1606
rect 2853 -1698 2860 -1523
rect 3024 -1608 3048 -1420
rect 3145 -1559 3158 -1369
rect 3240 -1423 3307 -1239
rect 3576 -1359 3723 697
rect 3573 -1427 3723 -1359
rect 3145 -1578 3157 -1559
rect 3210 -1578 3217 -1574
rect 3145 -1588 3218 -1578
rect 3210 -1598 3217 -1588
rect 3024 -1610 3155 -1608
rect 3024 -1624 3188 -1610
rect 3147 -1626 3188 -1624
rect 3179 -1698 3188 -1626
rect 3210 -1703 3215 -1598
rect 2153 -1887 2165 -1766
rect 2337 -1838 2468 -1832
rect 2777 -1886 2830 -1877
rect 2153 -1914 2163 -1887
rect 2777 -1915 2788 -1886
rect 2320 -2359 2362 -2334
<< m3contact >>
rect 398 1199 405 1204
rect -693 1092 -659 1106
rect -387 1095 -355 1109
rect -806 991 -789 1008
rect -458 990 -382 1011
rect -89 832 -73 851
rect -179 741 -150 761
rect -259 699 -241 712
rect 849 1139 857 1150
rect 402 1098 410 1103
rect 1142 1252 1156 1290
rect 820 1023 827 1028
rect 874 1023 879 1028
rect 852 1012 858 1017
rect 403 996 410 1003
rect 814 931 820 939
rect 857 921 862 927
rect 877 913 883 920
rect 399 903 407 908
rect 796 840 803 847
rect 874 840 879 846
rect 853 830 859 835
rect 405 805 411 811
rect 574 805 587 819
rect 402 699 411 705
rect 623 701 635 714
rect -265 513 -236 564
rect -179 549 -153 572
rect -92 542 -67 574
rect -21 441 -8 449
rect 1107 662 1115 672
rect 2396 612 2413 624
rect 400 594 407 600
rect 690 593 699 608
rect 1141 498 1151 505
rect 772 484 786 494
rect 1989 518 1997 527
rect 1566 493 1578 504
rect 154 441 165 447
rect 351 432 363 438
rect 1989 446 1996 457
rect 1565 422 1577 434
rect 2405 439 2413 446
rect -595 327 -573 338
rect -25 329 -8 335
rect 389 329 394 334
rect -671 233 -647 246
rect -52 233 -28 247
rect 414 230 422 236
rect 1285 281 1295 290
rect 1711 282 1720 292
rect 2093 290 2107 297
rect -795 158 -768 178
rect -54 157 -42 176
rect 415 128 420 133
rect 415 33 423 38
rect -123 -73 -105 -54
rect -35 -72 -17 -53
rect -252 -180 -231 -158
rect -29 -180 -9 -162
rect -352 -244 -325 -216
rect -24 -245 -9 -216
rect 413 -64 422 -58
rect 413 -164 418 -159
rect 414 -276 420 -271
rect 1 -416 17 -404
rect -603 -544 -575 -517
rect 173 -422 184 -410
rect -685 -712 -648 -681
rect -791 -757 -767 -744
rect 8 -755 19 -747
rect 1305 -29 1324 -18
rect 1071 -64 1089 -49
rect 2024 -262 2051 -256
rect 146 -543 151 -538
rect 425 -542 431 -537
rect 580 -541 591 -531
rect 377 -643 385 -635
rect 421 -643 429 -635
rect 586 -637 594 -631
rect 428 -740 434 -735
rect 558 -739 568 -734
rect 422 -835 427 -830
rect 565 -837 575 -832
rect 424 -921 429 -916
rect 434 -1043 439 -1036
rect 425 -1148 431 -1143
rect 3022 -1420 3050 -1397
rect 1448 -1564 1460 -1555
rect 474 -1636 484 -1617
rect 2153 -1561 2166 -1552
rect 1448 -1663 1460 -1652
rect 2153 -1675 2166 -1655
rect 1448 -1726 1460 -1719
rect 2153 -1766 2166 -1751
rect 2331 -1838 2337 -1831
rect 2830 -1886 2840 -1877
<< metal3 >>
rect -605 1202 -581 1206
rect -373 1203 398 1204
rect -562 1202 398 1203
rect -605 1199 398 1202
rect -605 1197 284 1199
rect -605 1196 -306 1197
rect -605 1195 -336 1196
rect -806 841 -789 991
rect -806 708 -787 841
rect -690 793 -660 1092
rect -605 844 -581 1195
rect 574 1139 849 1150
rect -7 1103 185 1104
rect -355 1102 334 1103
rect -355 1098 402 1102
rect -355 1097 -2 1098
rect 159 1097 366 1098
rect 574 1022 587 1139
rect 742 1024 807 1025
rect -382 1003 -171 1004
rect -30 1003 251 1004
rect -382 996 403 1003
rect -188 995 93 996
rect -88 907 399 908
rect -607 811 -581 844
rect -89 903 399 907
rect -89 851 -74 903
rect 574 819 586 1022
rect 623 1018 807 1024
rect 827 1023 874 1028
rect 623 1017 820 1018
rect 623 999 636 1017
rect 798 1012 852 1017
rect 623 853 635 999
rect 820 932 874 937
rect 815 925 857 927
rect 689 922 857 925
rect 689 917 821 922
rect 869 923 874 932
rect 869 920 883 923
rect -690 742 -653 793
rect -806 661 -785 708
rect -803 563 -785 661
rect -687 690 -653 742
rect -803 535 -783 563
rect -801 430 -783 535
rect -801 390 -782 430
rect -800 178 -782 390
rect -687 246 -651 690
rect -607 353 -583 811
rect -179 810 355 811
rect -179 805 405 810
rect -179 803 355 805
rect -179 761 -154 803
rect 623 714 634 853
rect 689 754 700 917
rect 803 840 874 846
rect 771 830 853 834
rect 771 759 786 830
rect -241 704 349 706
rect -241 699 402 704
rect 312 636 325 638
rect 312 630 406 636
rect 312 605 325 630
rect -364 594 325 605
rect 400 600 406 630
rect 690 608 699 754
rect -364 593 320 594
rect -607 338 -581 353
rect -607 327 -595 338
rect -687 233 -671 246
rect -800 158 -795 178
rect -800 37 -782 158
rect -800 16 -781 37
rect -799 -98 -781 16
rect -799 -136 -780 -98
rect -798 -349 -780 -136
rect -799 -393 -780 -349
rect -799 -485 -781 -393
rect -799 -522 -780 -485
rect -798 -592 -780 -522
rect -798 -652 -778 -592
rect -687 -609 -651 233
rect -607 169 -581 327
rect -605 75 -581 169
rect -605 -42 -579 75
rect -603 -517 -579 -42
rect -361 -216 -340 593
rect -265 -158 -241 513
rect -178 -54 -156 549
rect 771 562 785 759
rect 1142 735 1154 1252
rect 1141 701 1154 735
rect -91 452 -72 542
rect 772 494 785 562
rect 1107 672 1115 673
rect -91 431 -70 452
rect -8 441 154 447
rect 1107 438 1115 662
rect 1141 505 1151 701
rect 363 432 1121 438
rect 1566 434 1577 493
rect 1989 457 1996 518
rect 2405 446 2413 612
rect -90 133 -70 431
rect -8 329 389 333
rect 1071 290 1089 291
rect 1106 290 1296 291
rect 1550 290 1711 291
rect 1071 282 1285 290
rect 1071 279 1113 282
rect 1295 282 1296 290
rect 1432 289 1711 290
rect 1416 282 1711 289
rect 2092 290 2093 297
rect 1416 281 1589 282
rect -28 234 375 247
rect -28 233 414 234
rect 371 230 414 233
rect 1071 231 1089 279
rect 245 176 369 177
rect -42 157 369 176
rect -90 52 -68 133
rect 360 132 368 157
rect 360 128 415 132
rect -90 51 262 52
rect -90 39 377 51
rect -90 21 -68 39
rect 373 37 377 39
rect 373 33 415 37
rect -88 -36 -68 21
rect -178 -73 -123 -54
rect -178 -74 -106 -73
rect -265 -180 -252 -158
rect -361 -244 -352 -216
rect -798 -658 -776 -652
rect -796 -744 -776 -658
rect -685 -681 -651 -609
rect -796 -757 -791 -744
rect -796 -758 -776 -757
rect -361 -1144 -340 -244
rect -265 -1036 -241 -180
rect -178 -917 -156 -74
rect -88 -77 -66 -36
rect 1070 -49 1087 231
rect 1416 -19 1434 281
rect 2092 198 2107 290
rect 2048 195 2107 198
rect 1324 -29 1434 -19
rect 2024 184 2107 195
rect 2024 116 2053 184
rect 1306 -30 1433 -29
rect -17 -72 327 -54
rect -33 -74 327 -72
rect -88 -199 -68 -77
rect 312 -78 327 -74
rect 339 -64 413 -59
rect 1070 -60 1071 -49
rect 339 -65 374 -64
rect 339 -78 349 -65
rect 312 -83 349 -78
rect 321 -160 336 -159
rect 321 -163 413 -160
rect -9 -164 413 -163
rect -9 -179 336 -164
rect -9 -180 331 -179
rect -89 -424 -68 -199
rect -9 -245 364 -217
rect 358 -273 364 -245
rect 2024 -256 2051 116
rect 2024 -263 2051 -262
rect 358 -276 414 -273
rect 358 -278 364 -276
rect 17 -412 161 -404
rect 17 -416 173 -412
rect 151 -422 173 -416
rect -88 -494 -68 -424
rect -88 -684 -66 -494
rect 671 -531 1145 -530
rect 151 -542 425 -539
rect 671 -532 1174 -531
rect 591 -541 1174 -532
rect 151 -543 385 -542
rect 1061 -628 1076 -627
rect 728 -631 1076 -628
rect 385 -643 421 -635
rect 594 -636 1076 -631
rect 728 -637 1076 -636
rect -88 -853 -65 -684
rect 1061 -710 1076 -637
rect 970 -734 1002 -732
rect 361 -740 428 -736
rect 568 -739 1002 -734
rect 361 -748 370 -740
rect 19 -755 370 -748
rect -87 -874 -65 -853
rect 367 -835 422 -831
rect 367 -874 373 -835
rect 848 -833 868 -832
rect 714 -834 868 -833
rect 575 -837 868 -834
rect 714 -838 868 -837
rect -87 -888 373 -874
rect -178 -921 424 -917
rect -265 -1037 361 -1036
rect -265 -1043 434 -1037
rect 848 -1122 868 -838
rect 970 -1006 1002 -739
rect 1061 -900 1077 -710
rect 1147 -866 1174 -541
rect 1935 -856 2465 -853
rect 1757 -857 2465 -856
rect 1757 -860 2724 -857
rect 1589 -863 2724 -860
rect 1589 -865 3008 -863
rect 1299 -866 3008 -865
rect 1147 -889 3051 -866
rect 1147 -896 1568 -889
rect 2329 -892 3051 -889
rect 1062 -960 1077 -900
rect 3014 -905 3051 -892
rect 3022 -910 3051 -905
rect 1062 -963 1901 -960
rect 1062 -986 2842 -963
rect 970 -1009 1507 -1006
rect 970 -1014 1570 -1009
rect 2009 -1014 2024 -1009
rect 970 -1040 2024 -1014
rect 1033 -1043 2024 -1040
rect 848 -1123 1152 -1122
rect 848 -1124 1459 -1123
rect -361 -1145 -66 -1144
rect -361 -1148 425 -1145
rect 848 -1147 1460 -1124
rect 1096 -1148 1460 -1147
rect -361 -1149 -66 -1148
rect 1448 -1230 1460 -1148
rect 2009 -1213 2024 -1043
rect 2830 -1015 2840 -986
rect 2009 -1226 2166 -1213
rect 1448 -1309 1461 -1230
rect 2153 -1252 2166 -1226
rect 2830 -1246 2839 -1015
rect 3024 -1173 3046 -910
rect 3024 -1234 3047 -1173
rect 2153 -1262 2167 -1252
rect 2152 -1307 2167 -1262
rect 1448 -1519 1460 -1309
rect 2152 -1314 2166 -1307
rect 1448 -1555 1459 -1519
rect 2153 -1552 2166 -1314
rect 1867 -1614 2016 -1613
rect 997 -1615 1171 -1614
rect 1730 -1615 2016 -1614
rect 524 -1616 778 -1615
rect 839 -1616 1171 -1615
rect 1200 -1616 1502 -1615
rect 1730 -1616 2243 -1615
rect 524 -1617 2340 -1616
rect 484 -1635 2340 -1617
rect 484 -1636 1013 -1635
rect 1098 -1636 1879 -1635
rect 1992 -1636 2340 -1635
rect 2830 -1632 2840 -1246
rect 3024 -1397 3048 -1234
rect 691 -1637 865 -1636
rect 1098 -1637 1272 -1636
rect 1427 -1637 1757 -1636
rect 1448 -1719 1459 -1663
rect 2153 -1751 2165 -1675
rect 2331 -1789 2339 -1636
rect 2331 -1831 2337 -1789
rect 2830 -1877 2839 -1632
use decoder  decoder_0
timestamp 1699649695
transform 1 0 41 0 1 202
box -41 -202 165 271
use enable  enable_0
timestamp 1701060155
transform 0 1 406 -1 0 1265
box -28 -38 774 92
use enable  enable_1
timestamp 1701060155
transform 0 1 420 -1 0 396
box -28 -38 774 92
use enable  enable_2
timestamp 1701060155
transform 0 1 432 -1 0 -474
box -28 -38 774 92
use and_block  and_block_0
timestamp 1699691262
transform 0 1 843 -1 0 1073
box -27 -8 333 75
use 2_input_OR  2_input_OR_0
timestamp 1699680002
transform 1 0 101 0 1 -77
box -23 -24 68 39
use comparator_equal  comparator_equal_0
timestamp 1700304769
transform 1 0 1166 0 1 309
box -49 -1499 1958 182
use adder_subtractor  adder_subtractor_0
timestamp 1700257825
transform 1 0 3231 0 1 -1819
box -2047 -635 612 166
use 2_input_AND  2_input_AND_0
timestamp 1699478438
transform 1 0 3140 0 1 535
box -12 -30 69 33
<< labels >>
rlabel metal1 443 1373 455 1383 1 VDD
rlabel metal1 384 -1461 390 -1457 1 GND
rlabel metal1 888 739 890 740 1 AND_OUTPUT_A3B3
rlabel metal1 886 927 888 928 1 AND_OUTPUT_A1B1
rlabel metal1 886 1016 888 1017 1 AND_OUTPUT_A0B0
rlabel metal1 2878 -87 2880 -84 1 COMPARATOR_OUT_A_GREATERTHAN_B
rlabel metal1 2158 -1163 2160 -1160 1 COMPARATOR_OUT_A_LESSTHAN_B
rlabel metal1 27 220 29 222 1 S0_DECODER
rlabel metal1 170 262 172 264 1 S1_DECODER
rlabel metal1 109 484 110 485 1 S0_S1_DECODER
rlabel metal1 91 365 92 366 1 S0BAR_S1_DECODER
rlabel metal2 63 110 64 111 1 S0BAR_S1BAR_DECODER
rlabel metal1 113 -11 115 -10 1 S0_S1BAR_DECODER
rlabel metal1 396 1304 397 1305 1 INPUT_ALU_A0
rlabel metal3 346 1201 347 1202 1 INPUT_ALU_A1
rlabel metal3 351 1098 352 1099 1 INPUT_ALU_A2
rlabel metal3 353 999 354 1000 1 INPUT_ALU_A3
rlabel metal3 354 905 355 906 1 INPUT_ALU_B0
rlabel metal3 350 805 351 806 1 INPUT_ALU_B1
rlabel metal3 356 700 357 701 1 INPUT_ALU_B2
rlabel metal3 349 632 350 633 1 INPUT_ALU_B3
rlabel metal2 512 1201 513 1202 1 OUTPUT_ALU_ANDBLOCK_A0
rlabel metal2 513 1097 514 1098 1 OUTPUT_ALU_ANDBLOCK_A1
rlabel metal2 516 996 517 997 1 OUTPUT_ALU_ANDBLOCK_A2
rlabel metal2 519 902 520 903 1 OUTPUT_ALU_ANDBLOCK_A3
rlabel metal2 513 809 514 810 1 OUTPUT_ALU_ANDBLOCK_B0
rlabel metal2 519 704 520 705 1 OUTPUT_ALU_ANDBLOCK_B1
rlabel metal2 522 596 523 597 1 OUTPUT_ALU_ANDBLOCK_B2
rlabel metal2 524 487 525 488 1 OUTPUT_ALU_ANDBLOCK_B3
rlabel metal2 522 332 523 333 1 OUTPUT_ALU_COMPARATOR_A0
rlabel metal2 528 236 529 237 1 OUTPUT_ALU_COMPARATOR_A1
rlabel metal2 535 134 536 135 1 OUTPUT_ALU_COMPARATOR_A2
rlabel metal2 538 36 539 37 1 OUTPUT_ALU_COMPARATOR_A3
rlabel metal2 527 -59 528 -58 1 OUTPUT_ALU_COMPARATOR_B0
rlabel metal2 528 -164 529 -163 1 OUTPUT_ALU_COMPARATOR_B1
rlabel metal2 531 -268 532 -267 1 OUTPUT_ALU_COMPARATOR_B2
rlabel metal1 532 -380 533 -379 1 OUTPUT_ALU_COMPARATOR_B3
rlabel metal2 550 -536 551 -535 1 OUTPUT_ALU_ADDER_A0
rlabel metal2 559 -635 560 -634 1 OUTPUT_ALU_ADDER_A1
rlabel metal2 548 -738 549 -737 1 OUTPUT_ALU_ADDER_A2
rlabel metal2 549 -836 550 -835 1 OUTPUT_ALU_ADDER_A3
rlabel metal2 558 -930 559 -929 1 OUTPUT_ALU_ADDER_B0
rlabel metal2 552 -1034 553 -1033 1 OUTPUT_ALU_ADDER_B1
rlabel metal2 549 -1139 550 -1138 1 OUTPUT_ALU_ADDER_B2
rlabel metal2 476 -1275 477 -1274 1 OUTPUT_ALU_ADDER_B3
rlabel metal1 886 834 888 835 1 AND_OUTPUT_A2B2
rlabel m2contact 2888 403 2890 404 1 COMPARATOR_OUT_A_EQUAL_B
rlabel metal1 3216 536 3217 537 1 COMPARATOR_A_EQUAL_B_FINAL
rlabel metal1 3680 -1944 3683 -1942 1 ADDER_SUB_S0
rlabel metal1 3627 -1667 3634 -1665 1 ADD_SUB_M
rlabel metal1 3515 -2225 3517 -2223 1 ADDER_SUB_C1
rlabel metal1 3018 -1967 3020 -1966 1 ADDER_SUB_S1
rlabel metal1 2927 -2255 2930 -2253 1 ADDER_SUB_C2
rlabel metal1 2413 -1964 2414 -1963 1 ADDER_SUB_S2
rlabel metal1 2311 -2247 2313 -2246 1 ADDER_SUB_C3
rlabel metal1 1702 -1842 1704 -1840 1 ADDER_SUB_S3
rlabel metal1 1596 -2127 1599 -2125 1 ADDER_SUB_C4
rlabel metal1 1628 -2359 1630 -2357 1 ADDER_SUB_CFINAL
<< end >>
