* SPICE3 file created from enable.ext - technology: scmos
.include TSMC_180nm.txt


.param SUPPLY = 1.8


.global GND
.option scale=0.09u
Vdd VDD GND 'SUPPLY'
V_in_A0 A0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_A1 A1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
V_in_A2 A2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
V_in_A3 A3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)
V_in_enable enable gnd DC 0
* V_in_b0 node_b0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
* V_in_b1 node_b1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
* V_in_b2 node_b2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
* V_in_b3 node_b3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)

V_in_B0 B0 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_B1 B1 gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 140ns)
V_in_B2 B2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_B3 B3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)

M1000 VDD enable 2_input_AND_7/OUT 2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=672 pd=528 as=24 ps=20
M1001 2_input_AND_7/a_4_n21# B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=384 ps=320
M1002 B3_FINAL 2_input_AND_7/OUT VDD 2_input_AND_7/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1003 2_input_AND_7/OUT B3 VDD 2_input_AND_7/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 B3_FINAL 2_input_AND_7/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 2_input_AND_7/OUT enable 2_input_AND_7/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1006 VDD enable 2_input_AND_0/OUT 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1007 2_input_AND_0/a_4_n21# A0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1008 A0_FINAL 2_input_AND_0/OUT VDD 2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1009 2_input_AND_0/OUT A0 VDD 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 A0_FINAL 2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1011 2_input_AND_0/OUT enable 2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1012 VDD enable 2_input_AND_1/OUT 2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1013 2_input_AND_1/a_4_n21# A1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1014 A1_FINAL 2_input_AND_1/OUT VDD 2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1015 2_input_AND_1/OUT A1 VDD 2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 A1_FINAL 2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1017 2_input_AND_1/OUT enable 2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1018 VDD enable 2_input_AND_3/OUT 2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1019 2_input_AND_3/a_4_n21# A3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1020 A3_FINAL 2_input_AND_3/OUT VDD 2_input_AND_3/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1021 2_input_AND_3/OUT A3 VDD 2_input_AND_3/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 A3_FINAL 2_input_AND_3/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1023 2_input_AND_3/OUT enable 2_input_AND_3/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1024 VDD enable 2_input_AND_2/OUT 2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1025 2_input_AND_2/a_4_n21# A2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1026 A2_FINAL 2_input_AND_2/OUT VDD 2_input_AND_2/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1027 2_input_AND_2/OUT A2 VDD 2_input_AND_2/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 A2_FINAL 2_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1029 2_input_AND_2/OUT enable 2_input_AND_2/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1030 VDD enable 2_input_AND_4/OUT 2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1031 2_input_AND_4/a_4_n21# B0 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1032 B0_FINAL 2_input_AND_4/OUT VDD 2_input_AND_4/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1033 2_input_AND_4/OUT B0 VDD 2_input_AND_4/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 B0_FINAL 2_input_AND_4/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1035 2_input_AND_4/OUT enable 2_input_AND_4/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1036 VDD enable 2_input_AND_5/OUT 2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1037 2_input_AND_5/a_4_n21# B1 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1038 B1_FINAL 2_input_AND_5/OUT VDD 2_input_AND_5/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1039 2_input_AND_5/OUT B1 VDD 2_input_AND_5/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 B1_FINAL 2_input_AND_5/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1041 2_input_AND_5/OUT enable 2_input_AND_5/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1042 VDD enable 2_input_AND_6/OUT 2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1043 2_input_AND_6/a_4_n21# B2 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1044 B2_FINAL 2_input_AND_6/OUT VDD 2_input_AND_6/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1045 2_input_AND_6/OUT B2 VDD 2_input_AND_6/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 B2_FINAL 2_input_AND_6/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1047 2_input_AND_6/OUT enable 2_input_AND_6/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
C0 2_input_AND_5/OUT 2_input_AND_5/w_35_9# 0.08fF
C1 VDD A2_FINAL 0.02fF
C2 VDD 2_input_AND_3/OUT 0.06fF
C3 GND B2 0.05fF
C4 VDD 2_input_AND_0/OUT 0.06fF
C5 A0_FINAL 2_input_AND_0/w_35_9# 0.03fF
C6 2_input_AND_4/w_n12_9# enable 0.07fF
C7 2_input_AND_2/w_35_9# 2_input_AND_2/OUT 0.08fF
C8 GND A2 0.05fF
C9 GND 2_input_AND_4/OUT 0.04fF
C10 A1_FINAL 2_input_AND_1/w_35_9# 0.03fF
C11 2_input_AND_3/OUT 2_input_AND_3/w_n12_9# 0.03fF
C12 B1 enable 0.39fF
C13 2_input_AND_5/w_n12_9# enable 0.07fF
C14 VDD 2_input_AND_4/w_n12_9# 0.06fF
C15 2_input_AND_7/w_n12_9# 2_input_AND_7/OUT 0.03fF
C16 B2 2_input_AND_6/w_n12_9# 0.07fF
C17 GND 2_input_AND_6/OUT 0.04fF
C18 VDD 2_input_AND_5/w_n12_9# 0.06fF
C19 2_input_AND_1/OUT 2_input_AND_1/w_35_9# 0.08fF
C20 B2 enable 0.38fF
C21 GND B1_FINAL 0.05fF
C22 GND A0_FINAL 0.05fF
C23 2_input_AND_2/w_n12_9# A2 0.07fF
C24 B0_FINAL 2_input_AND_4/OUT 0.05fF
C25 GND 2_input_AND_7/OUT 0.04fF
C26 A2 enable 0.38fF
C27 2_input_AND_4/OUT enable 0.12fF
C28 VDD 2_input_AND_1/w_35_9# 0.03fF
C29 A0 2_input_AND_0/w_n12_9# 0.07fF
C30 2_input_AND_6/w_n12_9# 2_input_AND_6/OUT 0.03fF
C31 VDD 2_input_AND_4/OUT 0.06fF
C32 B3_FINAL 2_input_AND_7/OUT 0.05fF
C33 2_input_AND_6/OUT enable 0.12fF
C34 GND 2_input_AND_2/OUT 0.04fF
C35 GND A3 0.05fF
C36 GND A0 0.05fF
C37 VDD 2_input_AND_6/OUT 0.06fF
C38 2_input_AND_7/OUT enable 0.12fF
C39 2_input_AND_7/w_35_9# 2_input_AND_7/OUT 0.08fF
C40 GND A3_FINAL 0.05fF
C41 VDD B1_FINAL 0.02fF
C42 VDD A0_FINAL 0.02fF
C43 B2_FINAL 2_input_AND_6/OUT 0.05fF
C44 GND 2_input_AND_5/OUT 0.04fF
C45 B0_FINAL 2_input_AND_4/w_35_9# 0.03fF
C46 VDD 2_input_AND_7/OUT 0.06fF
C47 2_input_AND_5/w_n12_9# B1 0.07fF
C48 2_input_AND_2/w_n12_9# 2_input_AND_2/OUT 0.03fF
C49 VDD 2_input_AND_5/w_35_9# 0.03fF
C50 2_input_AND_2/OUT enable 0.12fF
C51 2_input_AND_3/w_35_9# A3_FINAL 0.03fF
C52 A3 enable 0.39fF
C53 GND B0 0.05fF
C54 A0 enable 0.38fF
C55 VDD 2_input_AND_4/w_35_9# 0.03fF
C56 VDD 2_input_AND_2/OUT 0.06fF
C57 2_input_AND_4/OUT 2_input_AND_4/w_n12_9# 0.03fF
C58 A0_FINAL 2_input_AND_0/OUT 0.05fF
C59 2_input_AND_5/OUT enable 0.12fF
C60 B3 2_input_AND_7/w_n12_9# 0.07fF
C61 A3 2_input_AND_3/w_n12_9# 0.07fF
C62 VDD A3_FINAL 0.02fF
C63 VDD 2_input_AND_5/OUT 0.06fF
C64 A1 2_input_AND_1/w_n12_9# 0.07fF
C65 B0 enable 0.39fF
C66 VDD 2_input_AND_2/w_35_9# 0.03fF
C67 VDD 2_input_AND_6/w_35_9# 0.03fF
C68 A2_FINAL 2_input_AND_2/OUT 0.05fF
C69 A1 GND 0.05fF
C70 GND B3 0.05fF
C71 B2_FINAL 2_input_AND_6/w_35_9# 0.03fF
C72 2_input_AND_7/w_n12_9# enable 0.07fF
C73 VDD 2_input_AND_0/w_35_9# 0.03fF
C74 GND A1_FINAL 0.05fF
C75 enable 2_input_AND_0/w_n12_9# 0.07fF
C76 GND B3_FINAL 0.05fF
C77 A3_FINAL 2_input_AND_3/OUT 0.05fF
C78 2_input_AND_1/OUT 2_input_AND_1/w_n12_9# 0.03fF
C79 2_input_AND_2/w_35_9# A2_FINAL 0.03fF
C80 2_input_AND_1/w_n12_9# enable 0.07fF
C81 VDD 2_input_AND_7/w_n12_9# 0.07fF
C82 VDD 2_input_AND_0/w_n12_9# 0.06fF
C83 GND B0_FINAL 0.05fF
C84 GND 2_input_AND_1/OUT 0.04fF
C85 A1 enable 0.39fF
C86 GND enable 3.23fF
C87 VDD 2_input_AND_1/w_n12_9# 0.06fF
C88 B3 enable 0.41fF
C89 2_input_AND_1/OUT A1_FINAL 0.05fF
C90 2_input_AND_0/w_35_9# 2_input_AND_0/OUT 0.08fF
C91 2_input_AND_4/OUT 2_input_AND_4/w_35_9# 0.08fF
C92 2_input_AND_5/w_n12_9# 2_input_AND_5/OUT 0.03fF
C93 2_input_AND_7/w_35_9# B3_FINAL 0.03fF
C94 B0 2_input_AND_4/w_n12_9# 0.07fF
C95 GND B2_FINAL 0.05fF
C96 2_input_AND_2/w_n12_9# enable 0.07fF
C97 VDD A1_FINAL 0.02fF
C98 VDD 2_input_AND_3/w_35_9# 0.03fF
C99 2_input_AND_6/w_n12_9# enable 0.07fF
C100 VDD B3_FINAL 0.02fF
C101 2_input_AND_1/OUT enable 0.12fF
C102 2_input_AND_0/OUT 2_input_AND_0/w_n12_9# 0.03fF
C103 2_input_AND_5/w_35_9# B1_FINAL 0.03fF
C104 2_input_AND_2/w_n12_9# VDD 0.06fF
C105 VDD 2_input_AND_6/w_n12_9# 0.07fF
C106 VDD B0_FINAL 0.02fF
C107 GND A2_FINAL 0.05fF
C108 VDD 2_input_AND_1/OUT 0.06fF
C109 GND 2_input_AND_3/OUT 0.04fF
C110 GND 2_input_AND_0/OUT 0.04fF
C111 VDD 2_input_AND_7/w_35_9# 0.03fF
C112 2_input_AND_3/w_n12_9# enable 0.07fF
C113 2_input_AND_3/w_35_9# 2_input_AND_3/OUT 0.08fF
C114 2_input_AND_6/OUT 2_input_AND_6/w_35_9# 0.08fF
C115 VDD B2_FINAL 0.02fF
C116 VDD 2_input_AND_3/w_n12_9# 0.06fF
C117 GND B1 0.05fF
C118 2_input_AND_5/OUT B1_FINAL 0.05fF
C119 2_input_AND_3/OUT enable 0.12fF
C120 2_input_AND_0/OUT enable 0.12fF
C121 GND Gnd 8.47fF
C122 VDD Gnd 5.85fF
C123 B2_FINAL Gnd 0.12fF
C124 2_input_AND_6/OUT Gnd 0.38fF
C125 B2 Gnd 0.26fF
C126 2_input_AND_6/w_35_9# Gnd 0.56fF
C127 2_input_AND_6/w_n12_9# Gnd 0.72fF
C128 B1_FINAL Gnd 0.12fF
C129 2_input_AND_5/OUT Gnd 0.38fF
C130 B1 Gnd 0.22fF
C131 2_input_AND_5/w_35_9# Gnd 0.56fF
C132 2_input_AND_5/w_n12_9# Gnd 0.72fF
C133 B0_FINAL Gnd 0.12fF
C134 2_input_AND_4/OUT Gnd 0.38fF
C135 B0 Gnd 0.22fF
C136 2_input_AND_4/w_35_9# Gnd 0.56fF
C137 2_input_AND_4/w_n12_9# Gnd 0.72fF
C138 A2_FINAL Gnd 0.12fF
C139 2_input_AND_2/OUT Gnd 0.38fF
C140 A2 Gnd 0.25fF
C141 2_input_AND_2/w_35_9# Gnd 0.56fF
C142 2_input_AND_2/w_n12_9# Gnd 0.72fF
C143 A3_FINAL Gnd 0.11fF
C144 2_input_AND_3/OUT Gnd 0.38fF
C145 A3 Gnd 0.25fF
C146 2_input_AND_3/w_35_9# Gnd 0.56fF
C147 2_input_AND_3/w_n12_9# Gnd 0.72fF
C148 A1_FINAL Gnd 0.12fF
C149 2_input_AND_1/OUT Gnd 0.38fF
C150 A1 Gnd 0.25fF
C151 2_input_AND_1/w_35_9# Gnd 0.56fF
C152 2_input_AND_1/w_n12_9# Gnd 0.72fF
C153 A0_FINAL Gnd 0.12fF
C154 2_input_AND_0/OUT Gnd 0.38fF
C155 enable Gnd 2.47fF
C156 A0 Gnd 0.25fF
C157 2_input_AND_0/w_35_9# Gnd 0.56fF
C158 2_input_AND_0/w_n12_9# Gnd 0.72fF
C159 B3_FINAL Gnd 0.10fF
C160 2_input_AND_7/OUT Gnd 0.38fF
C161 B3 Gnd 0.26fF
C162 2_input_AND_7/w_35_9# Gnd 0.56fF
C163 2_input_AND_7/w_n12_9# Gnd 0.72fF
.tran 1n 500n
.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6 
plot v(B0) v(B1)+2 v(B2)+4 v(B3)+6
plot v(A0_FINAL) v(A1_FINAL)+2 v(A2_FINAL)+4 v(A3_FINAL)+6 
plot v(B0_FINAL) v(B1_FINAL)+2 v(B2_FINAL)+4 v(B3_FINAL)+6
* plot v(A0_BAR_A1_BAR) v(A0_A1_BAR)+2 v(A0_BAR_A1)+4 v(A0_A1)+6
* plot v(OUT_FINAL)/
* hardcopy image.ps v(node_a) v(node_b)+2 v(OUT)+4
.end
.endc