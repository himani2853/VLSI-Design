magic
tech scmos
timestamp 1699649695
<< metal1 >>
rect 46 267 62 271
rect 46 265 50 267
rect 53 177 57 196
rect -8 172 57 177
rect 60 178 64 196
rect 60 172 127 178
rect -8 30 -2 172
rect 48 157 62 161
rect 48 155 52 157
rect 55 71 59 85
rect 41 66 59 71
rect 62 71 66 84
rect 122 71 127 172
rect 62 66 127 71
rect 41 30 46 66
rect 122 34 127 66
rect -8 26 7 30
rect 28 26 46 30
rect -8 -97 -2 26
rect 22 4 27 10
rect 22 -14 28 4
rect 41 -4 46 26
rect 73 30 93 34
rect 112 30 127 34
rect 73 -3 78 30
rect 41 -8 54 -4
rect 22 -18 39 -14
rect 50 -23 54 -8
rect 57 -8 120 -3
rect 57 -22 61 -8
rect 56 -93 68 -90
rect 115 -97 120 -8
rect -8 -102 58 -97
rect 54 -116 58 -102
rect 61 -102 120 -97
rect 61 -116 65 -102
rect 63 -188 72 -184
<< m2contact >>
rect 17 185 22 191
rect 75 185 80 192
rect 72 121 77 126
rect 19 75 24 80
rect 5 50 11 56
rect 88 50 95 56
rect 109 50 114 56
rect 27 4 34 10
rect 101 4 107 9
rect 92 -23 98 -18
rect 97 -110 102 -105
rect 42 -183 48 -176
<< metal2 >>
rect -26 185 17 188
rect -26 181 22 185
rect 80 185 165 188
rect 75 182 165 185
rect -26 56 -16 181
rect 150 126 165 182
rect 77 121 165 126
rect 5 75 19 80
rect 5 56 11 75
rect 150 56 165 121
rect -41 50 5 56
rect 50 50 88 56
rect 114 50 165 56
rect -41 49 -16 50
rect 50 49 95 50
rect -41 5 -26 49
rect 50 10 58 49
rect -40 -2 -26 5
rect 34 4 58 10
rect 101 -2 107 4
rect -40 -9 107 -2
rect 101 -18 107 -9
rect 98 -23 107 -18
rect 102 -110 107 -23
rect 150 -108 165 50
rect 43 -192 48 -183
rect 149 -192 164 -108
rect 43 -202 164 -192
use q1a_NOT  q1a_NOT_0
timestamp 1698924755
transform 1 0 17 0 1 27
box -12 -23 15 29
use q1a_NOT  q1a_NOT_1
timestamp 1698924755
transform -1 0 103 0 -1 33
box -12 -23 15 29
use 2_input_AND  2_input_AND_0
timestamp 1699478438
transform 0 1 64 -1 0 -23
box -12 -30 69 33
use 2_input_AND  2_input_AND_1
timestamp 1699478438
transform 0 1 68 -1 0 -117
box -12 -30 69 33
use 2_input_AND  2_input_AND_2
timestamp 1699478438
transform 0 -1 52 1 0 87
box -12 -30 69 33
use 2_input_AND  2_input_AND_3
timestamp 1699478438
transform 0 -1 50 1 0 197
box -12 -30 69 33
<< labels >>
rlabel metal1 -6 27 -5 28 1 A0
rlabel metal1 124 32 125 33 1 A1
rlabel metal1 75 19 76 20 1 A1_BAR
rlabel metal1 42 28 43 29 1 A0_BAR
rlabel metal2 -35 31 -34 32 1 VDD
rlabel metal2 159 37 160 38 1 GND
rlabel metal1 61 -92 61 -92 1 A0_BAR_A1_BAR
rlabel metal1 55 159 56 160 1 A0_BAR_A1
rlabel metal1 67 -187 68 -186 1 A0_A1_BAR
rlabel metal1 55 268 56 269 5 A0_A1
<< end >>
