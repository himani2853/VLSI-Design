magic
tech scmos
timestamp 1699478438
<< nwell >>
rect -12 9 28 27
rect 35 9 69 27
<< ntransistor >>
rect 52 -13 54 -9
rect 2 -21 4 -17
rect 10 -21 12 -17
<< ptransistor >>
rect 2 16 4 20
rect 10 16 12 20
rect 52 16 54 20
<< ndiffusion >>
rect 50 -13 52 -9
rect 54 -13 56 -9
rect 0 -21 2 -17
rect 4 -21 10 -17
rect 12 -21 16 -17
<< pdiffusion >>
rect 0 16 2 20
rect 4 16 5 20
rect 9 16 10 20
rect 12 16 16 20
rect 49 16 52 20
rect 54 16 56 20
<< ndcontact >>
rect 46 -13 50 -9
rect 56 -13 60 -9
rect -4 -21 0 -17
rect 16 -21 20 -17
<< pdcontact >>
rect -4 16 0 20
rect 5 16 9 20
rect 16 16 20 20
rect 45 16 49 20
rect 56 16 60 20
<< polysilicon >>
rect 2 20 4 23
rect 10 20 12 23
rect 52 20 54 24
rect 2 -3 4 16
rect 2 -17 4 -7
rect 10 -10 12 16
rect 52 4 54 16
rect 53 0 54 4
rect 52 -9 54 0
rect 10 -17 12 -14
rect 52 -16 54 -13
rect 2 -27 4 -21
rect 10 -27 12 -21
<< polycontact >>
rect 0 -7 4 -3
rect 48 0 53 4
rect 8 -14 12 -10
<< metal1 >>
rect -12 28 69 33
rect -4 20 0 28
rect 16 20 20 28
rect 45 20 49 28
rect 5 4 9 16
rect 56 4 60 16
rect 5 0 48 4
rect 56 0 69 4
rect -3 -7 0 -3
rect -3 -14 8 -10
rect 16 -17 20 0
rect 56 -9 60 0
rect 46 -20 50 -13
rect -4 -25 0 -21
rect 28 -25 66 -20
rect -11 -30 33 -25
<< labels >>
rlabel metal1 33 30 34 31 5 VDD
rlabel metal1 -1 -5 0 -4 1 A
rlabel metal1 0 -12 1 -11 1 B
rlabel metal1 37 1 38 2 1 OUT
rlabel metal1 65 2 66 3 7 OUT_FINAL
rlabel metal1 24 -29 25 -28 1 GND
<< end >>
