* SPICE3 file created from comparator_equal.ext - technology: scmos
.include TSMC_180nm.txt


.param SUPPLY = 1.8


.global GND

Vdd VDD GND 'SUPPLY'
V_in_A0 A0 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_B0 B0 GND PULSE(0 1.8 0ns 100ps 100ps 100ns 200ns)
V_in_A1 A1 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_B1 B1 GND PULSE(0 1.8 0ns 100ps 100ps 100ns 200ns)
V_in_A2 A2 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_B2 B2 GND PULSE(0 1.8 0ns 100ps 100ps 100ns 200ns)
V_in_A3 A3 GND PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_B3 B3 GND PULSE(0 1.8 0ns 100ps 100ps 100ns 200ns)
* V_in_A0 A0 GND DC 1.8
* V_in_A1 A1 GND DC 0
* V_in_A2 A2 GND DC 0
* V_in_A3 A3 GND DC 1.8

* V_in_B0 B0 GND DC 1.8
* V_in_B1 B1 GND DC 1.8
* V_in_B2 B2 GND DC 1.8
* V_in_B3 B3 GND DC 1.8

.option scale=0.09u

M1000 B0_NOT B0 VDD q1a_NOT_3/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=2058 ps=1258
M1001 B0_NOT B0 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=1965 ps=1146
M1002 q1a_NOT_4/out A3 VDD q1a_NOT_4/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1003 q1a_NOT_4/out A3 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1004 A2NOT q1a_NOT_5/in VDD q1a_NOT_5/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1005 A2NOT q1a_NOT_5/in GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1006 A0NOT A0 VDD q1a_NOT_6/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1007 A0NOT A0 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1008 A1NOT A1 VDD q1a_NOT_7/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1009 A1NOT A1 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1010 VDD A2B2 q1b_5_INPUT_AND_0/OUT q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=154 ps=86
M1011 q1b_5_INPUT_AND_0/OUT A0 VDD q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 q1b_5_INPUT_AND_0/OUT A1B1 VDD q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1b_5_INPUT_AND_0/OUT GND Gnd CMOSN w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1014 q1b_5_INPUT_AND_0/a_n11_n43# A3B3 GND Gnd CMOSN w=7 l=2
+  ad=56 pd=30 as=0 ps=0
M1015 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1b_5_INPUT_AND_0/OUT VDD q1b_5_INPUT_AND_0/w_50_10# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1016 q1b_5_INPUT_AND_0/a_n1_n43# A2B2 q1b_5_INPUT_AND_0/a_n11_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1017 q1b_5_INPUT_AND_0/OUT A0 q1b_5_INPUT_AND_0/a_17_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1018 q1b_5_INPUT_AND_0/a_17_n43# B0_NOT q1b_5_INPUT_AND_0/a_8_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1019 q1b_5_INPUT_AND_0/OUT A3B3 VDD q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 VDD B0_NOT q1b_5_INPUT_AND_0/OUT q1b_5_INPUT_AND_0/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 q1b_5_INPUT_AND_0/a_8_n43# A1B1 q1b_5_INPUT_AND_0/a_n1_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 VDD A2B2 q1b_5_INPUT_AND_1/OUT q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=154 ps=86
M1023 q1b_5_INPUT_AND_1/OUT A0NOT VDD q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1024 q1b_5_INPUT_AND_1/OUT A1B1 VDD q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 q1b_5_INPUT_AND_1/OUT GND Gnd CMOSN w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1026 q1b_5_INPUT_AND_1/a_n11_n43# A3B3 GND Gnd CMOSN w=7 l=2
+  ad=56 pd=30 as=0 ps=0
M1027 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 q1b_5_INPUT_AND_1/OUT VDD q1b_5_INPUT_AND_1/w_50_10# CMOSP w=6 l=2
+  ad=48 pd=28 as=0 ps=0
M1028 q1b_5_INPUT_AND_1/a_n1_n43# A2B2 q1b_5_INPUT_AND_1/a_n11_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1029 q1b_5_INPUT_AND_1/OUT A0NOT q1b_5_INPUT_AND_1/a_17_n43# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1030 q1b_5_INPUT_AND_1/a_17_n43# B0 q1b_5_INPUT_AND_1/a_8_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1031 q1b_5_INPUT_AND_1/OUT A3B3 VDD q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 VDD B0 q1b_5_INPUT_AND_1/OUT q1b_5_INPUT_AND_1/w_n24_8# CMOSP w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1033 q1b_5_INPUT_AND_1/a_8_n43# A1B1 q1b_5_INPUT_AND_1/a_n1_n43# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 A_greater_than_B q1c_4_INPUT_OR_0/OUT VDD q1c_4_INPUT_OR_0/w_41_n9# CMOSP w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1035 GND A3_B3NOT q1c_4_INPUT_OR_0/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=270 ps=114
M1036 q1c_4_INPUT_OR_0/OUT A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1c_4_INPUT_OR_0/a_1_0# q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=90 pd=38 as=90 ps=38
M1037 q1c_4_INPUT_OR_0/OUT A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 q1c_4_INPUT_OR_0/OUT A2_B2NOT_A3B3XNOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 q1c_4_INPUT_OR_0/a_n18_0# A3_B3NOT VDD q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1040 q1c_4_INPUT_OR_0/a_1_0# A1_B1NOT_A3B3XNOR_A2B2XOR q1c_4_INPUT_OR_0/a_n9_0# q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1041 A_greater_than_B q1c_4_INPUT_OR_0/OUT GND Gnd CMOSN w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1042 q1c_4_INPUT_OR_0/a_n9_0# A2_B2NOT_A3B3XNOR q1c_4_INPUT_OR_0/a_n18_0# q1c_4_INPUT_OR_0/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 GND A1_B1NOT_A3B3XNOR_A2B2XOR q1c_4_INPUT_OR_0/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 A_less_than_B q1c_4_INPUT_OR_1/OUT VDD q1c_4_INPUT_OR_1/w_41_n9# CMOSP w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1045 GND A3NOT_B3 q1c_4_INPUT_OR_1/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=270 ps=114
M1046 q1c_4_INPUT_OR_1/OUT A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 q1c_4_INPUT_OR_1/a_1_0# q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=90 pd=38 as=90 ps=38
M1047 q1c_4_INPUT_OR_1/OUT A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 q1c_4_INPUT_OR_1/OUT A2NOT_B2_A3B3XNOR GND Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1049 q1c_4_INPUT_OR_1/a_n18_0# A3NOT_B3 VDD q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 q1c_4_INPUT_OR_1/a_1_0# A1NOTB1_A2XNORB2_A3XNORB3 q1c_4_INPUT_OR_1/a_n9_0# q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=80 ps=36
M1051 A_less_than_B q1c_4_INPUT_OR_1/OUT GND Gnd CMOSN w=8 l=3
+  ad=112 pd=44 as=0 ps=0
M1052 q1c_4_INPUT_OR_1/a_n9_0# A2NOT_B2_A3B3XNOR q1c_4_INPUT_OR_1/a_n18_0# q1c_4_INPUT_OR_1/w_n38_n10# CMOSP w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 GND A1NOTB1_A2XNORB2_A3XNORB3 q1c_4_INPUT_OR_1/OUT Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 4_input_AND_0/a_n8_n45# A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1055 4_input_AND_0/OUT A2B2 VDD 4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=0 ps=0
M1056 A_IS_EQUAL_B 4_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1057 VDD A3B3 4_input_AND_0/OUT 4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 4_input_AND_0/OUT A0B0 4_input_AND_0/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1059 VDD A1B1 4_input_AND_0/OUT 4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 A_IS_EQUAL_B 4_input_AND_0/OUT VDD 4_input_AND_0/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1061 4_input_AND_0/a_10_n45# A1B1 4_input_AND_0/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1062 4_input_AND_0/OUT A0B0 VDD 4_input_AND_0/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 4_input_AND_0/a_1_n45# A2B2 4_input_AND_0/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 3_input_AND_0/OUT A2 3_input_AND_0/a_6_n34# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=24 ps=20
M1065 3_input_AND_0/OUT A2 VDD 3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=56 pd=44 as=0 ps=0
M1066 3_input_AND_0/a_6_n34# B2_NOT 3_input_AND_0/a_n3_n34# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=28 ps=22
M1067 VDD B2_NOT 3_input_AND_0/OUT 3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 3_input_AND_0/OUT A3B3 VDD 3_input_AND_0/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 A2_B2NOT_A3B3XNOR 3_input_AND_0/OUT VDD 3_input_AND_0/w_34_3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1070 A2_B2NOT_A3B3XNOR 3_input_AND_0/OUT GND Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1071 3_input_AND_0/a_n3_n34# A3B3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 4_input_AND_1/a_n8_n45# A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1073 4_input_AND_1/OUT A2B2 q1a_NOT_2/vdd 4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=142 ps=96
M1074 A1_B1NOT_A3B3XNOR_A2B2XOR 4_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1075 q1a_NOT_2/vdd A3B3 4_input_AND_1/OUT 4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1076 4_input_AND_1/OUT A1 4_input_AND_1/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1077 q1a_NOT_2/vdd B1_NOT 4_input_AND_1/OUT 4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 A1_B1NOT_A3B3XNOR_A2B2XOR 4_input_AND_1/OUT q1a_NOT_2/vdd 4_input_AND_1/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1079 4_input_AND_1/a_10_n45# B1_NOT 4_input_AND_1/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1080 4_input_AND_1/OUT A1 q1a_NOT_2/vdd 4_input_AND_1/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 4_input_AND_1/a_1_n45# A2B2 4_input_AND_1/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 VDD B1 XNOR_1/q1d_2_INPUT_XOR_0/BBAR XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1083 XNOR_1/OUT XNOR_1/q1d_2_INPUT_XOR_0/BBAR XNOR_1/q1d_2_INPUT_XOR_0/ABAR XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1084 XNOR_1/q1d_2_INPUT_XOR_0/BBAR B1 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1085 VDD A1 XNOR_1/q1d_2_INPUT_XOR_0/ABAR XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 XNOR_1/OUT B1 A1 XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=24 ps=20
M1087 XNOR_1/q1d_2_INPUT_XOR_0/ABAR A1 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1088 XNOR_1/OUT XNOR_1/q1d_2_INPUT_XOR_0/BBAR A1 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=24 ps=20
M1089 XNOR_1/OUT B1 XNOR_1/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1090 A1B1 XNOR_1/OUT VDD XNOR_1/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1091 A1B1 XNOR_1/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1092 VDD B0 XNOR_0/q1d_2_INPUT_XOR_0/BBAR XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1093 XNOR_0/OUT XNOR_0/q1d_2_INPUT_XOR_0/BBAR XNOR_0/q1d_2_INPUT_XOR_0/ABAR XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1094 XNOR_0/q1d_2_INPUT_XOR_0/BBAR B0 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1095 VDD A0 XNOR_0/q1d_2_INPUT_XOR_0/ABAR XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 XNOR_0/OUT B0 A0 XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=24 ps=20
M1097 XNOR_0/q1d_2_INPUT_XOR_0/ABAR A0 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1098 XNOR_0/OUT XNOR_0/q1d_2_INPUT_XOR_0/BBAR A0 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=24 ps=20
M1099 XNOR_0/OUT B0 XNOR_0/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1100 A0B0 XNOR_0/OUT VDD XNOR_0/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1101 A0B0 XNOR_0/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1102 VDD A3 2_input_AND_0/OUT 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1103 2_input_AND_0/a_4_n21# B3_NOT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1104 A3_B3NOT 2_input_AND_0/OUT VDD 2_input_AND_0/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1105 2_input_AND_0/OUT B3_NOT VDD 2_input_AND_0/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 A3_B3NOT 2_input_AND_0/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1107 2_input_AND_0/OUT A3 2_input_AND_0/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1108 3_input_AND_1/OUT A2NOT 3_input_AND_1/a_6_n34# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=24 ps=20
M1109 3_input_AND_1/OUT A2NOT VDD 3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=56 pd=44 as=0 ps=0
M1110 3_input_AND_1/a_6_n34# B2 3_input_AND_1/a_n3_n34# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=28 ps=22
M1111 VDD B2 3_input_AND_1/OUT 3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 3_input_AND_1/OUT A3B3 VDD 3_input_AND_1/w_n19_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 A2NOT_B2_A3B3XNOR 3_input_AND_1/OUT VDD 3_input_AND_1/w_34_3# CMOSP w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1114 A2NOT_B2_A3B3XNOR 3_input_AND_1/OUT GND Gnd CMOSN w=5 l=2
+  ad=30 pd=22 as=0 ps=0
M1115 3_input_AND_1/a_n3_n34# A3B3 GND Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 4_input_AND_2/a_n8_n45# A3B3 GND Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=0 ps=0
M1117 4_input_AND_2/OUT A2B2 VDD 4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=102 pd=70 as=0 ps=0
M1118 A1NOTB1_A2XNORB2_A3XNORB3 4_input_AND_2/OUT GND Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1119 VDD A3B3 4_input_AND_2/OUT 4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 4_input_AND_2/OUT A1NOT 4_input_AND_2/a_10_n45# Gnd CMOSN w=7 l=2
+  ad=49 pd=28 as=49 ps=28
M1121 VDD B1 4_input_AND_2/OUT 4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 A1NOTB1_A2XNORB2_A3XNORB3 4_input_AND_2/OUT VDD 4_input_AND_2/w_40_5# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1123 4_input_AND_2/a_10_n45# B1 4_input_AND_2/a_1_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=49 ps=28
M1124 4_input_AND_2/OUT A1NOT VDD 4_input_AND_2/w_n22_4# CMOSP w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 4_input_AND_2/a_1_n45# A2B2 4_input_AND_2/a_n8_n45# Gnd CMOSN w=7 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 VDD B2 XNOR_2/q1d_2_INPUT_XOR_0/BBAR XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1127 XNOR_2/OUT XNOR_2/q1d_2_INPUT_XOR_0/BBAR XNOR_2/q1d_2_INPUT_XOR_0/ABAR XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1128 XNOR_2/q1d_2_INPUT_XOR_0/BBAR B2 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1129 VDD A2 XNOR_2/q1d_2_INPUT_XOR_0/ABAR XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 XNOR_2/OUT B2 A2 XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=24 ps=20
M1131 XNOR_2/q1d_2_INPUT_XOR_0/ABAR A2 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1132 XNOR_2/OUT XNOR_2/q1d_2_INPUT_XOR_0/BBAR A2 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=24 ps=20
M1133 XNOR_2/OUT B2 XNOR_2/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1134 A2B2 XNOR_2/OUT VDD XNOR_2/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1135 A2B2 XNOR_2/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1136 VDD q1a_NOT_4/out 2_input_AND_1/OUT 2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1137 2_input_AND_1/a_4_n21# B3 GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1138 A3NOT_B3 2_input_AND_1/OUT VDD 2_input_AND_1/w_35_9# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1139 2_input_AND_1/OUT B3 VDD 2_input_AND_1/w_n12_9# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 A3NOT_B3 2_input_AND_1/OUT GND Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1141 2_input_AND_1/OUT q1a_NOT_4/out 2_input_AND_1/a_4_n21# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1142 VDD B3 XNOR_3/q1d_2_INPUT_XOR_0/BBAR XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1143 XNOR_3/OUT XNOR_3/q1d_2_INPUT_XOR_0/BBAR XNOR_3/q1d_2_INPUT_XOR_0/ABAR XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# CMOSP w=4 l=3
+  ad=52 pd=42 as=44 ps=38
M1144 XNOR_3/q1d_2_INPUT_XOR_0/BBAR B3 GND Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1145 VDD A3 XNOR_3/q1d_2_INPUT_XOR_0/ABAR XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 XNOR_3/OUT B3 A3 XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# CMOSP w=4 l=3
+  ad=0 pd=0 as=24 ps=20
M1147 XNOR_3/q1d_2_INPUT_XOR_0/ABAR A3 GND Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=0 ps=0
M1148 XNOR_3/OUT XNOR_3/q1d_2_INPUT_XOR_0/BBAR A3 Gnd CMOSN w=4 l=3
+  ad=48 pd=40 as=24 ps=20
M1149 XNOR_3/OUT B3 XNOR_3/q1d_2_INPUT_XOR_0/ABAR Gnd CMOSN w=4 l=3
+  ad=0 pd=0 as=0 ps=0
M1150 A3B3 XNOR_3/OUT VDD XNOR_3/w_181_105# CMOSP w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1151 A3B3 XNOR_3/OUT GND Gnd CMOSN w=7 l=4
+  ad=126 pd=50 as=0 ps=0
M1152 B3_NOT B3 VDD q1a_NOT_0/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1153 B3_NOT B3 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1154 B2_NOT B2 VDD q1a_NOT_1/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1155 B2_NOT B2 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1156 B1_NOT B1 q1a_NOT_2/vdd q1a_NOT_2/w_n12_4# CMOSP w=6 l=2
+  ad=36 pd=24 as=0 ps=0
M1157 B1_NOT B1 GND Gnd CMOSN w=6 l=2
+  ad=36 pd=24 as=0 ps=0
C0 A1B1 B1 0.32fF
C1 q1a_NOT_5/in A2NOT 0.04fF
C2 VDD 4_input_AND_0/w_n22_4# 0.05fF
C3 q1a_NOT_2/vdd 4_input_AND_1/w_n22_4# 0.05fF
C4 4_input_AND_1/OUT 4_input_AND_1/w_40_5# 0.07fF
C5 XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# B3 0.09fF
C6 3_input_AND_1/w_n19_2# A3B3 0.08fF
C7 VDD q1c_4_INPUT_OR_0/w_n38_n10# 0.11fF
C8 XNOR_1/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C9 q1a_NOT_2/vdd B1_NOT 0.10fF
C10 A2 GND 0.75fF
C11 VDD B1 0.45fF
C12 A3B3 A2_B2NOT_A3B3XNOR 0.75fF
C13 XNOR_0/q1d_2_INPUT_XOR_0/ABAR XNOR_0/OUT 0.19fF
C14 A0 GND 0.20fF
C15 VDD XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C16 A1NOTB1_A2XNORB2_A3XNORB3 A3B3 0.30fF
C17 q1a_NOT_5/in GND 0.04fF
C18 q1c_4_INPUT_OR_1/w_n38_n10# q1c_4_INPUT_OR_1/OUT 0.06fF
C19 A2 q1a_NOT_5/in 0.72fF
C20 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1b_5_INPUT_AND_0/OUT 0.05fF
C21 XNOR_3/OUT XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C22 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A1 0.19fF
C23 B3_NOT 2_input_AND_0/w_n12_9# 0.07fF
C24 2_input_AND_0/OUT A3_B3NOT 0.05fF
C25 XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C26 VDD 3_input_AND_0/OUT 0.09fF
C27 A1NOT A2B2 0.08fF
C28 XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# XNOR_2/OUT 0.03fF
C29 A3NOT_B3 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C30 XNOR_2/OUT XNOR_2/w_181_105# 0.13fF
C31 A0B0 B3 0.19fF
C32 B1 GND 0.87fF
C33 XNOR_1/q1d_2_INPUT_XOR_0/BBAR B1 0.03fF
C34 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A1B1 0.33fF
C35 A1_B1NOT_A3B3XNOR_A2B2XOR B3 0.17fF
C36 4_input_AND_2/OUT A1NOT 0.14fF
C37 XNOR_0/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C38 XNOR_1/q1d_2_INPUT_XOR_0/ABAR XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C39 A3NOT_B3 2_input_AND_1/w_35_9# 0.03fF
C40 XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# B3 0.08fF
C41 A_greater_than_B GND 0.05fF
C42 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR VDD 0.07fF
C43 A2NOT_B2_A3B3XNOR 3_input_AND_1/OUT 0.05fF
C44 VDD A3NOT_B3 0.02fF
C45 q1c_4_INPUT_OR_1/w_41_n9# A_less_than_B 0.05fF
C46 GND 3_input_AND_0/OUT 0.09fF
C47 VDD XNOR_2/w_181_105# 0.06fF
C48 XNOR_0/w_181_105# XNOR_0/OUT 0.13fF
C49 A3B3 A2B2 5.18fF
C50 4_input_AND_0/w_40_5# 4_input_AND_0/OUT 0.07fF
C51 A1NOTB1_A2XNORB2_A3XNORB3 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 1.40fF
C52 A2 3_input_AND_0/OUT 0.13fF
C53 q1c_4_INPUT_OR_0/OUT A3_B3NOT 0.09fF
C54 3_input_AND_0/w_n19_2# B2_NOT 0.08fF
C55 B0 XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# 0.09fF
C56 3_input_AND_0/w_34_3# VDD 0.03fF
C57 B2_NOT q1a_NOT_1/w_n12_4# 0.04fF
C58 XNOR_2/OUT XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C59 B0 A3B3 0.08fF
C60 B0 q1a_NOT_3/w_n12_4# 0.09fF
C61 VDD XNOR_3/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C62 A0B0 4_input_AND_0/OUT 0.14fF
C63 VDD 2_input_AND_0/w_n12_9# 0.06fF
C64 3_input_AND_1/w_34_3# 3_input_AND_1/OUT 0.06fF
C65 VDD 3_input_AND_1/w_n19_2# 0.06fF
C66 XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C67 4_input_AND_2/OUT A3B3 0.15fF
C68 XNOR_3/q1d_2_INPUT_XOR_0/ABAR XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# 0.03fF
C69 B2_NOT A3B3 0.50fF
C70 VDD A2_B2NOT_A3B3XNOR 0.06fF
C71 VDD 2_input_AND_0/w_35_9# 0.03fF
C72 3_input_AND_1/w_n19_2# A2NOT 0.08fF
C73 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR GND 0.14fF
C74 B0_NOT A3B3 0.08fF
C75 A1NOTB1_A2XNORB2_A3XNORB3 4_input_AND_2/w_40_5# 0.03fF
C76 q1a_NOT_3/w_n12_4# B0_NOT 0.04fF
C77 A3NOT_B3 GND 0.11fF
C78 q1a_NOT_2/vdd A3B3 0.12fF
C79 q1a_NOT_4/out 2_input_AND_1/w_n12_9# 0.07fF
C80 VDD XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C81 q1c_4_INPUT_OR_1/w_n38_n10# A2NOT_B2_A3B3XNOR 0.10fF
C82 XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# A2 0.03fF
C83 A0B0 XNOR_0/w_181_105# 0.06fF
C84 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1a_NOT_5/in 0.21fF
C85 A1_B1NOT_A3B3XNOR_A2B2XOR A3_B3NOT 0.09fF
C86 A1 4_input_AND_1/a_1_n45# 0.01fF
C87 XNOR_3/q1d_2_INPUT_XOR_0/ABAR GND 0.23fF
C88 q1b_5_INPUT_AND_0/OUT A2B2 0.17fF
C89 A1 A2B2 0.34fF
C90 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1b_5_INPUT_AND_0/w_50_10# 0.04fF
C91 XNOR_3/w_181_105# A3B3 0.06fF
C92 XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# VDD 0.03fF
C93 XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# XNOR_0/OUT 0.03fF
C94 A_less_than_B GND 0.04fF
C95 A0NOT A3B3 0.08fF
C96 4_input_AND_1/w_n22_4# B1_NOT 0.08fF
C97 GND A2_B2NOT_A3B3XNOR 0.10fF
C98 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1c_4_INPUT_OR_0/w_n38_n10# 0.10fF
C99 XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C100 B2 q1a_NOT_1/w_n12_4# 0.10fF
C101 q1a_NOT_4/out VDD 0.46fF
C102 A3B3 A3 0.29fF
C103 A1NOT 4_input_AND_2/w_n22_4# 0.07fF
C104 A1NOTB1_A2XNORB2_A3XNORB3 GND 0.06fF
C105 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR B1 0.16fF
C106 A1B1 A2B2 4.95fF
C107 XNOR_2/q1d_2_INPUT_XOR_0/ABAR GND 0.23fF
C108 B2 A3B3 3.41fF
C109 q1b_5_INPUT_AND_0/OUT B0_NOT 0.08fF
C110 B3 A3_B3NOT 0.15fF
C111 A2 XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C112 A1 XNOR_1/OUT 0.18fF
C113 A1B1 B0 1.08fF
C114 XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.09fF
C115 XNOR_3/OUT XNOR_3/w_181_105# 0.13fF
C116 XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# XNOR_3/OUT 0.03fF
C117 VDD A2B2 1.39fF
C118 q1b_5_INPUT_AND_1/w_n24_8# A3B3 0.09fF
C119 q1c_4_INPUT_OR_1/OUT A2NOT_B2_A3B3XNOR 0.09fF
C120 XNOR_2/q1d_2_INPUT_XOR_0/BBAR B2 0.03fF
C121 B0 VDD 0.27fF
C122 VDD q1a_NOT_4/w_n12_4# 0.08fF
C123 XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# A2 0.08fF
C124 XNOR_3/OUT A3 0.18fF
C125 q1c_4_INPUT_OR_0/w_n38_n10# A2_B2NOT_A3B3XNOR 0.10fF
C126 B3_NOT A3 0.57fF
C127 A0B0 A3B3 0.34fF
C128 XNOR_0/q1d_2_INPUT_XOR_0/ABAR XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C129 4_input_AND_1/OUT A2B2 0.09fF
C130 4_input_AND_2/OUT 4_input_AND_2/w_40_5# 0.07fF
C131 XNOR_3/q1d_2_INPUT_XOR_0/BBAR XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C132 VDD 4_input_AND_2/OUT 0.21fF
C133 q1a_NOT_4/out GND 0.50fF
C134 XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# A3 0.08fF
C135 A3B3 4_input_AND_2/w_n22_4# 0.28fF
C136 A1B1 B0_NOT 0.73fF
C137 XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_2/OUT 0.04fF
C138 VDD XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C139 A1_B1NOT_A3B3XNOR_A2B2XOR A3B3 1.07fF
C140 VDD B2_NOT 0.10fF
C141 VDD 2_input_AND_0/OUT 0.06fF
C142 q1b_5_INPUT_AND_1/OUT A2B2 0.17fF
C143 A1 XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C144 3_input_AND_0/w_34_3# 3_input_AND_0/OUT 0.06fF
C145 VDD B0_NOT 0.10fF
C146 q1b_5_INPUT_AND_1/OUT B0 0.08fF
C147 2_input_AND_1/w_n12_9# 2_input_AND_1/OUT 0.03fF
C148 VDD 3_input_AND_1/OUT 0.09fF
C149 A2B2 GND 1.52fF
C150 XNOR_3/q1d_2_INPUT_XOR_0/BBAR B3 0.03fF
C151 A2_B2NOT_A3B3XNOR 3_input_AND_0/OUT 0.05fF
C152 A0 A2B2 0.08fF
C153 B0 GND 1.36fF
C154 4_input_AND_1/OUT q1a_NOT_2/vdd 0.21fF
C155 A0NOT A1B1 0.08fF
C156 A0NOT q1a_NOT_6/w_n12_4# 0.09fF
C157 2_input_AND_1/OUT 2_input_AND_1/w_35_9# 0.08fF
C158 XNOR_2/OUT B2 0.15fF
C159 A2NOT 3_input_AND_1/OUT 0.13fF
C160 A1B1 A3 0.17fF
C161 B0 A0 0.43fF
C162 q1a_NOT_5/in A2B2 0.31fF
C163 4_input_AND_2/OUT GND 0.11fF
C164 q1c_4_INPUT_OR_1/w_n38_n10# A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C165 q1b_5_INPUT_AND_0/w_n24_8# A3B3 0.09fF
C166 XNOR_3/w_181_105# VDD 0.06fF
C167 A3B3 B3 0.22fF
C168 B2_NOT GND 0.12fF
C169 VDD XNOR_0/OUT 0.17fF
C170 VDD 2_input_AND_1/OUT 0.06fF
C171 VDD XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C172 2_input_AND_0/OUT GND 0.04fF
C173 A0NOT VDD 0.10fF
C174 B2_NOT A2 0.38fF
C175 A1 A0B0 0.38fF
C176 A1B1 B2 0.18fF
C177 VDD A3 0.01fF
C178 B0_NOT GND 0.10fF
C179 4_input_AND_0/w_n22_4# A2B2 0.07fF
C180 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A2_B2NOT_A3B3XNOR 0.10fF
C181 A0 B0_NOT 0.84fF
C182 3_input_AND_1/OUT GND 0.09fF
C183 4_input_AND_1/w_n22_4# A3B3 0.07fF
C184 A1B1 q1b_5_INPUT_AND_1/w_n24_8# 0.07fF
C185 VDD B2 0.81fF
C186 B1 A2B2 2.42fF
C187 q1c_4_INPUT_OR_1/w_n38_n10# VDD 0.11fF
C188 A3B3 B1_NOT 0.08fF
C189 A3NOT_B3 A1NOTB1_A2XNORB2_A3XNORB3 0.09fF
C190 A0NOT q1b_5_INPUT_AND_1/OUT 0.13fF
C191 A1B1 A0B0 1.20fF
C192 XNOR_3/OUT B3 0.15fF
C193 B3_NOT B3 0.04fF
C194 XNOR_1/OUT XNOR_1/w_181_105# 0.13fF
C195 3_input_AND_0/w_34_3# A2_B2NOT_A3B3XNOR 0.03fF
C196 VDD q1b_5_INPUT_AND_1/w_n24_8# 0.15fF
C197 VDD 4_input_AND_0/w_40_5# 0.03fF
C198 q1a_NOT_2/vdd 4_input_AND_1/w_40_5# 0.03fF
C199 q1a_NOT_2/w_n12_4# B1 0.10fF
C200 A2NOT B2 0.39fF
C201 4_input_AND_0/OUT A3B3 0.15fF
C202 VDD q1c_4_INPUT_OR_0/w_41_n9# 0.09fF
C203 A1_B1NOT_A3B3XNOR_A2B2XOR A1B1 0.58fF
C204 4_input_AND_2/OUT B1 0.09fF
C205 B0 XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C206 2_input_AND_1/OUT GND 0.04fF
C207 XNOR_1/q1d_2_INPUT_XOR_0/ABAR GND 0.23fF
C208 A1 XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C209 A0NOT GND 0.27fF
C210 VDD A0B0 0.42fF
C211 VDD 4_input_AND_2/w_n22_4# 0.05fF
C212 q1b_5_INPUT_AND_0/w_n24_8# q1b_5_INPUT_AND_0/OUT 0.08fF
C213 A3 GND 0.79fF
C214 A0 XNOR_0/OUT 0.18fF
C215 XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# B2 0.08fF
C216 q1c_4_INPUT_OR_0/OUT GND 0.63fF
C217 A0NOT A0 0.04fF
C218 XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# XNOR_0/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C219 q1c_4_INPUT_OR_1/OUT A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.78fF
C220 XNOR_1/OUT B1 0.15fF
C221 q1b_5_INPUT_AND_1/OUT q1b_5_INPUT_AND_1/w_n24_8# 0.08fF
C222 VDD XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C223 2_input_AND_1/w_n12_9# B3 0.07fF
C224 q1c_4_INPUT_OR_1/w_41_n9# q1c_4_INPUT_OR_1/OUT 0.10fF
C225 B2 GND 1.19fF
C226 3_input_AND_1/w_34_3# A2NOT_B2_A3B3XNOR 0.03fF
C227 A2 B2 0.30fF
C228 A1_B1NOT_A3B3XNOR_A2B2XOR 4_input_AND_1/OUT 0.04fF
C229 q1b_5_INPUT_AND_1/w_50_10# A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.04fF
C230 A3B3 A3_B3NOT 0.15fF
C231 A1 4_input_AND_1/w_n22_4# 0.07fF
C232 B2_NOT 3_input_AND_0/OUT 0.08fF
C233 A1B1 q1b_5_INPUT_AND_0/w_n24_8# 0.07fF
C234 A1B1 B3 0.19fF
C235 XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_0/OUT 0.04fF
C236 A1 B1_NOT 0.37fF
C237 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A2B2 0.19fF
C238 A0B0 GND 1.64fF
C239 A2NOT_B2_A3B3XNOR A3B3 0.29fF
C240 XNOR_1/q1d_2_INPUT_XOR_0/ABAR B1 0.08fF
C241 q1c_4_INPUT_OR_0/OUT q1c_4_INPUT_OR_0/w_n38_n10# 0.06fF
C242 q1a_NOT_7/w_n12_4# A1NOT 0.04fF
C243 A2 A0B0 0.26fF
C244 VDD q1b_5_INPUT_AND_0/w_n24_8# 0.15fF
C245 VDD B3 1.46fF
C246 A1_B1NOT_A3B3XNOR_A2B2XOR GND 0.06fF
C247 XNOR_2/w_181_105# A2B2 0.06fF
C248 A1NOT A3B3 0.05fF
C249 VDD q1b_5_INPUT_AND_1/w_50_10# 0.06fF
C250 VDD XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C251 XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C252 A1 XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C253 A1_B1NOT_A3B3XNOR_A2B2XOR q1a_NOT_5/in 0.40fF
C254 A1_B1NOT_A3B3XNOR_A2B2XOR 4_input_AND_1/w_40_5# 0.03fF
C255 3_input_AND_0/w_n19_2# A3B3 0.08fF
C256 A1B1 4_input_AND_0/OUT 0.09fF
C257 4_input_AND_0/w_n22_4# A0B0 0.07fF
C258 A2B2 A2_B2NOT_A3B3XNOR 0.29fF
C259 q1b_5_INPUT_AND_1/OUT q1b_5_INPUT_AND_1/w_50_10# 0.07fF
C260 q1c_4_INPUT_OR_1/OUT GND 0.63fF
C261 4_input_AND_1/OUT 4_input_AND_1/w_n22_4# 0.09fF
C262 A1NOTB1_A2XNORB2_A3XNORB3 A2B2 0.25fF
C263 2_input_AND_0/w_n12_9# 2_input_AND_0/OUT 0.03fF
C264 A0B0 B1 0.15fF
C265 B3 GND 0.95fF
C266 A1_B1NOT_A3B3XNOR_A2B2XOR q1c_4_INPUT_OR_0/w_n38_n10# 0.10fF
C267 VDD 4_input_AND_0/OUT 0.21fF
C268 4_input_AND_1/OUT B1_NOT 0.09fF
C269 B1 4_input_AND_2/w_n22_4# 0.08fF
C270 XNOR_0/q1d_2_INPUT_XOR_0/ABAR GND 0.23fF
C271 q1b_5_INPUT_AND_0/w_n24_8# A0 0.07fF
C272 q1a_NOT_0/w_n12_4# B3 0.10fF
C273 A_greater_than_B q1c_4_INPUT_OR_0/w_41_n9# 0.05fF
C274 A1NOTB1_A2XNORB2_A3XNORB3 4_input_AND_2/OUT 0.04fF
C275 VDD XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C276 A0 XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C277 3_input_AND_1/w_n19_2# 3_input_AND_1/OUT 0.06fF
C278 2_input_AND_0/w_35_9# 2_input_AND_0/OUT 0.08fF
C279 2_input_AND_1/OUT A3NOT_B3 0.05fF
C280 A1 A1NOT 0.04fF
C281 A2NOT_B2_A3B3XNOR A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.10fF
C282 4_input_AND_0/w_40_5# A_IS_EQUAL_B 0.03fF
C283 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A3 0.47fF
C284 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR q1c_4_INPUT_OR_0/OUT 0.78fF
C285 VDD A3_B3NOT 0.02fF
C286 B1_NOT GND 0.23fF
C287 VDD XNOR_0/w_181_105# 0.06fF
C288 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR B2 0.26fF
C289 B1 XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# 0.09fF
C290 A2 3_input_AND_0/a_n3_n34# 0.01fF
C291 q1a_NOT_4/out q1a_NOT_4/w_n12_4# 0.04fF
C292 4_input_AND_0/OUT GND 0.11fF
C293 XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# B2 0.09fF
C294 XNOR_0/q1d_2_INPUT_XOR_0/ABAR XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# 0.03fF
C295 XNOR_3/q1d_2_INPUT_XOR_0/ABAR A3 0.08fF
C296 q1c_4_INPUT_OR_1/w_n38_n10# A3NOT_B3 0.13fF
C297 2_input_AND_0/w_n12_9# A3 0.07fF
C298 XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_1/OUT 0.04fF
C299 VDD XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.03fF
C300 VDD A2NOT_B2_A3B3XNOR 0.31fF
C301 q1a_NOT_7/w_n12_4# A1 0.12fF
C302 XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_2/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C303 q1b_5_INPUT_AND_0/OUT A3B3 0.05fF
C304 A1 A3B3 0.53fF
C305 VDD A1NOT 0.10fF
C306 A3 A2_B2NOT_A3B3XNOR 0.35fF
C307 3_input_AND_1/w_n19_2# B2 0.08fF
C308 q1c_4_INPUT_OR_0/OUT A2_B2NOT_A3B3XNOR 0.09fF
C309 B0 A2B2 0.08fF
C310 A1_B1NOT_A3B3XNOR_A2B2XOR A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR 1.20fF
C311 GND A3_B3NOT 0.11fF
C312 VDD 3_input_AND_1/w_34_3# 0.03fF
C313 4_input_AND_2/OUT A2B2 0.09fF
C314 B1 B1_NOT 0.04fF
C315 4_input_AND_0/w_n22_4# 4_input_AND_0/OUT 0.09fF
C316 XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.03fF
C317 3_input_AND_0/w_n19_2# VDD 0.06fF
C318 VDD q1a_NOT_1/w_n12_4# 0.07fF
C319 q1c_4_INPUT_OR_1/w_n38_n10# A1NOTB1_A2XNORB2_A3XNORB3 0.10fF
C320 A1B1 A3B3 1.84fF
C321 B0 XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# 0.08fF
C322 VDD XNOR_3/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C323 XNOR_2/q1d_2_INPUT_XOR_0/ABAR B2 0.08fF
C324 B0_NOT A2B2 0.08fF
C325 VDD q1a_NOT_7/w_n12_4# 0.07fF
C326 A2NOT_B2_A3B3XNOR GND 0.10fF
C327 q1a_NOT_2/vdd A2B2 0.11fF
C328 A0 XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# 0.08fF
C329 XNOR_3/q1d_2_INPUT_XOR_0/BBAR XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# 0.09fF
C330 B0 B0_NOT 0.04fF
C331 q1a_NOT_4/out 2_input_AND_1/OUT 0.12fF
C332 VDD A3B3 2.00fF
C333 VDD q1a_NOT_3/w_n12_4# 0.07fF
C334 A1NOT GND 0.13fF
C335 q1c_4_INPUT_OR_1/OUT A3NOT_B3 0.09fF
C336 q1a_NOT_4/out A3 0.04fF
C337 A1_B1NOT_A3B3XNOR_A2B2XOR A2_B2NOT_A3B3XNOR 1.54fF
C338 q1a_NOT_2/vdd q1a_NOT_2/w_n12_4# 0.05fF
C339 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR B3 0.63fF
C340 q1c_4_INPUT_OR_0/w_n38_n10# A3_B3NOT 0.12fF
C341 4_input_AND_1/OUT A3B3 0.15fF
C342 A2NOT A3B3 0.01fF
C343 VDD XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C344 4_input_AND_0/OUT A_IS_EQUAL_B 0.04fF
C345 q1b_5_INPUT_AND_1/OUT A3B3 0.05fF
C346 A0NOT A2B2 0.08fF
C347 VDD XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# 0.03fF
C348 XNOR_3/q1d_2_INPUT_XOR_0/ABAR B3 0.08fF
C349 XNOR_3/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C350 3_input_AND_0/w_n19_2# A2 0.08fF
C351 A2B2 A3 0.16fF
C352 B0 XNOR_0/OUT 0.15fF
C353 A0NOT B0 1.29fF
C354 XNOR_3/OUT VDD 0.12fF
C355 VDD B3_NOT 0.10fF
C356 q1a_NOT_4/w_n12_4# A3 0.09fF
C357 A1B1 q1b_5_INPUT_AND_0/OUT 0.08fF
C358 XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# VDD 0.03fF
C359 A3B3 GND 0.83fF
C360 A1B1 A1 0.36fF
C361 B2 A2B2 0.37fF
C362 XNOR_3/OUT XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# 0.04fF
C363 B3 A2_B2NOT_A3B3XNOR 0.18fF
C364 A0 XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C365 q1c_4_INPUT_OR_1/OUT A1NOTB1_A2XNORB2_A3XNORB3 0.17fF
C366 XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# XNOR_2/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C367 B1 A1NOT 0.67fF
C368 A0 A3B3 0.08fF
C369 VDD q1b_5_INPUT_AND_0/OUT 0.32fF
C370 A3 2_input_AND_0/OUT 0.12fF
C371 XNOR_1/OUT XNOR_1/q1d_2_INPUT_XOR_0/ABAR 0.19fF
C372 VDD A1 0.42fF
C373 q1b_5_INPUT_AND_1/w_n24_8# A2B2 0.07fF
C374 q1a_NOT_5/in A3B3 1.07fF
C375 XNOR_2/q1d_2_INPUT_XOR_0/BBAR GND 0.04fF
C376 XNOR_2/OUT VDD 0.13fF
C377 VDD 2_input_AND_1/w_n12_9# 0.06fF
C378 B0 q1b_5_INPUT_AND_1/w_n24_8# 0.07fF
C379 B2_NOT B2 0.04fF
C380 VDD A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.07fF
C381 A0B0 A2B2 0.35fF
C382 A1 4_input_AND_1/OUT 0.14fF
C383 XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C384 q1c_4_INPUT_OR_1/w_41_n9# VDD 0.20fF
C385 A2B2 4_input_AND_2/w_n22_4# 0.07fF
C386 A1_B1NOT_A3B3XNOR_A2B2XOR A2B2 0.74fF
C387 4_input_AND_0/w_n22_4# A3B3 0.07fF
C388 B3_NOT GND 0.15fF
C389 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A3_B3NOT 0.10fF
C390 A1B1 VDD 1.48fF
C391 VDD q1a_NOT_6/w_n12_4# 0.05fF
C392 VDD 2_input_AND_1/w_35_9# 0.03fF
C393 3_input_AND_1/OUT B2 0.08fF
C394 q1a_NOT_0/w_n12_4# B3_NOT 0.04fF
C395 B1 A3B3 0.54fF
C396 4_input_AND_2/OUT 4_input_AND_2/w_n22_4# 0.09fF
C397 q1a_NOT_4/out B3 1.40fF
C398 q1b_5_INPUT_AND_1/OUT A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 0.05fF
C399 VDD q1a_NOT_5/w_n12_4# 0.08fF
C400 XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# A3 0.03fF
C401 VDD 4_input_AND_2/w_40_5# 0.03fF
C402 q1b_5_INPUT_AND_0/OUT GND 0.06fF
C403 A1 GND 1.28fF
C404 3_input_AND_0/w_n19_2# 3_input_AND_0/OUT 0.06fF
C405 q1b_5_INPUT_AND_0/OUT A0 0.13fF
C406 A3NOT_B3 A2NOT_B2_A3B3XNOR 2.38fF
C407 q1b_5_INPUT_AND_1/OUT A1B1 0.08fF
C408 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 GND 0.14fF
C409 q1a_NOT_5/w_n12_4# A2NOT 0.04fF
C410 XNOR_2/OUT A2 0.18fF
C411 VDD A2NOT 0.10fF
C412 q1b_5_INPUT_AND_0/w_n24_8# A2B2 0.07fF
C413 A2B2 B3 0.28fF
C414 XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# B1 0.08fF
C415 A3_B3NOT A2_B2NOT_A3B3XNOR 2.07fF
C416 q1b_5_INPUT_AND_1/OUT VDD 0.32fF
C417 q1b_5_INPUT_AND_0/OUT q1b_5_INPUT_AND_0/w_50_10# 0.07fF
C418 2_input_AND_0/w_35_9# A3_B3NOT 0.03fF
C419 A1B1 GND 1.87fF
C420 A0NOT q1b_5_INPUT_AND_1/w_n24_8# 0.07fF
C421 XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# VDD 0.03fF
C422 A1B1 A2 0.27fF
C423 B0 XNOR_0/q1d_2_INPUT_XOR_0/ABAR 0.08fF
C424 q1a_NOT_6/w_n12_4# A0 0.09fF
C425 A1B1 A0 0.08fF
C426 q1c_4_INPUT_OR_0/OUT q1c_4_INPUT_OR_0/w_41_n9# 0.10fF
C427 XNOR_1/OUT XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# 0.03fF
C428 4_input_AND_1/w_n22_4# A2B2 0.07fF
C429 VDD GND 4.35fF
C430 VDD XNOR_1/q1d_2_INPUT_XOR_0/BBAR 0.03fF
C431 A0B0 A3 0.17fF
C432 VDD A2 0.01fF
C433 A1 B1 0.17fF
C434 VDD A0 0.01fF
C435 A2B2 B1_NOT 1.02fF
C436 A2NOT_B2_A3B3XNOR A1NOTB1_A2XNORB2_A3XNORB3 2.05fF
C437 q1b_5_INPUT_AND_0/w_n24_8# B0_NOT 0.07fF
C438 q1a_NOT_0/w_n12_4# VDD 0.07fF
C439 A1B1 XNOR_1/w_181_105# 0.06fF
C440 A1_B1NOT_A3B3XNOR_A2B2XOR A3 0.42fF
C441 q1a_NOT_5/w_n12_4# q1a_NOT_5/in 0.12fF
C442 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR A3B3 0.22fF
C443 A1_B1NOT_A3B3XNOR_A2B2XOR q1c_4_INPUT_OR_0/OUT 0.17fF
C444 4_input_AND_1/OUT GND 0.11fF
C445 B2 A0B0 0.18fF
C446 VDD q1a_NOT_5/in 0.44fF
C447 A2NOT GND 0.47fF
C448 4_input_AND_0/OUT A2B2 0.09fF
C449 A1B1 4_input_AND_0/w_n22_4# 0.08fF
C450 q1a_NOT_2/w_n12_4# B1_NOT 0.04fF
C451 VDD XNOR_1/w_181_105# 0.06fF
C452 A1_B1NOT_A3B3XNOR_A2B2XOR B2 0.48fF
C453 q1b_5_INPUT_AND_1/OUT GND 0.06fF
C454 VDD q1b_5_INPUT_AND_0/w_50_10# 0.06fF
C455 GND Gnd 68.11fF
C456 VDD Gnd 114.89fF
C457 q1a_NOT_2/w_n12_4# Gnd 0.50fF
C458 q1a_NOT_1/w_n12_4# Gnd 0.50fF
C459 q1a_NOT_0/w_n12_4# Gnd 0.50fF
C460 XNOR_3/w_181_105# Gnd 2.32fF
C461 XNOR_3/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C462 XNOR_3/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C463 XNOR_3/OUT Gnd 1.20fF
C464 XNOR_3/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C465 XNOR_3/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C466 XNOR_3/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C467 XNOR_3/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C468 2_input_AND_1/OUT Gnd 0.38fF
C469 q1a_NOT_4/out Gnd 0.58fF
C470 B3 Gnd 2.34fF
C471 2_input_AND_1/w_35_9# Gnd 0.56fF
C472 2_input_AND_1/w_n12_9# Gnd 0.72fF
C473 XNOR_2/w_181_105# Gnd 2.32fF
C474 XNOR_2/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C475 XNOR_2/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C476 XNOR_2/OUT Gnd 1.20fF
C477 A2 Gnd 7.85fF
C478 XNOR_2/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C479 XNOR_2/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C480 XNOR_2/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C481 XNOR_2/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C482 4_input_AND_2/OUT Gnd 0.72fF
C483 A1NOT Gnd 0.93fF
C484 B1 Gnd 1.47fF
C485 A2B2 Gnd 2.49fF
C486 A3B3 Gnd 3.25fF
C487 4_input_AND_2/w_40_5# Gnd 0.51fF
C488 4_input_AND_2/w_n22_4# Gnd 0.99fF
C489 3_input_AND_1/OUT Gnd 0.51fF
C490 A2NOT Gnd 0.94fF
C491 B2 Gnd 1.38fF
C492 3_input_AND_1/w_34_3# Gnd 0.48fF
C493 3_input_AND_1/w_n19_2# Gnd 0.83fF
C494 2_input_AND_0/OUT Gnd 0.38fF
C495 B3_NOT Gnd 0.41fF
C496 2_input_AND_0/w_35_9# Gnd 0.56fF
C497 2_input_AND_0/w_n12_9# Gnd 0.72fF
C498 A0B0 Gnd 1.50fF
C499 XNOR_0/w_181_105# Gnd 2.32fF
C500 XNOR_0/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C501 XNOR_0/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C502 XNOR_0/OUT Gnd 1.20fF
C503 XNOR_0/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C504 XNOR_0/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C505 XNOR_0/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C506 XNOR_0/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C507 XNOR_1/w_181_105# Gnd 2.32fF
C508 XNOR_1/q1d_2_INPUT_XOR_0/ABAR Gnd 0.10fF
C509 XNOR_1/q1d_2_INPUT_XOR_0/BBAR Gnd 0.04fF
C510 XNOR_1/OUT Gnd 1.20fF
C511 XNOR_1/q1d_2_INPUT_XOR_0/w_53_n17# Gnd 0.45fF
C512 XNOR_1/q1d_2_INPUT_XOR_0/w_12_2# Gnd 0.04fF
C513 XNOR_1/q1d_2_INPUT_XOR_0/w_n34_1# Gnd 0.08fF
C514 XNOR_1/q1d_2_INPUT_XOR_0/w_52_34# Gnd 0.45fF
C515 q1a_NOT_2/vdd Gnd 0.59fF
C516 4_input_AND_1/OUT Gnd 0.72fF
C517 B1_NOT Gnd 0.67fF
C518 4_input_AND_1/w_40_5# Gnd 0.51fF
C519 4_input_AND_1/w_n22_4# Gnd 0.99fF
C520 3_input_AND_0/OUT Gnd 0.51fF
C521 B2_NOT Gnd 0.41fF
C522 3_input_AND_0/w_34_3# Gnd 0.48fF
C523 3_input_AND_0/w_n19_2# Gnd 0.83fF
C524 A_IS_EQUAL_B Gnd 0.10fF
C525 4_input_AND_0/OUT Gnd 0.72fF
C526 4_input_AND_0/w_40_5# Gnd 0.51fF
C527 4_input_AND_0/w_n22_4# Gnd 0.99fF
C528 A_less_than_B Gnd 0.26fF
C529 q1c_4_INPUT_OR_1/OUT Gnd 0.92fF
C530 A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3 Gnd 7.27fF
C531 A2NOT_B2_A3B3XNOR Gnd 4.26fF
C532 A3NOT_B3 Gnd 4.30fF
C533 q1c_4_INPUT_OR_1/w_41_n9# Gnd 1.25fF
C534 q1c_4_INPUT_OR_1/w_n38_n10# Gnd 1.97fF
C535 A_greater_than_B Gnd 0.33fF
C536 q1c_4_INPUT_OR_0/OUT Gnd 0.92fF
C537 A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR Gnd 13.09fF
C538 A1_B1NOT_A3B3XNOR_A2B2XOR Gnd 16.15fF
C539 A2_B2NOT_A3B3XNOR Gnd 7.25fF
C540 A3_B3NOT Gnd 1.55fF
C541 q1c_4_INPUT_OR_0/w_41_n9# Gnd 1.25fF
C542 q1c_4_INPUT_OR_0/w_n38_n10# Gnd 1.97fF
C543 q1b_5_INPUT_AND_1/OUT Gnd 0.31fF
C544 A0NOT Gnd 0.71fF
C545 B0 Gnd 1.67fF
C546 A1B1 Gnd 1.91fF
C547 q1b_5_INPUT_AND_1/w_50_10# Gnd 0.06fF
C548 q1b_5_INPUT_AND_1/w_n24_8# Gnd 1.35fF
C549 q1b_5_INPUT_AND_0/OUT Gnd 0.31fF
C550 B0_NOT Gnd 0.42fF
C551 q1b_5_INPUT_AND_0/w_50_10# Gnd 0.06fF
C552 q1b_5_INPUT_AND_0/w_n24_8# Gnd 1.35fF
C553 A1 Gnd 10.34fF
C554 q1a_NOT_7/w_n12_4# Gnd 0.50fF
C555 A0 Gnd 15.26fF
C556 q1a_NOT_6/w_n12_4# Gnd 0.50fF
C557 q1a_NOT_5/in Gnd 0.49fF
C558 q1a_NOT_5/w_n12_4# Gnd 0.50fF
C559 A3 Gnd 4.06fF
C560 q1a_NOT_4/w_n12_4# Gnd 0.50fF
C561 q1a_NOT_3/w_n12_4# Gnd 0.50fF
.tran 1n 500n

.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(A0) v(A1)+2 v(A2)+4 v(A3)+6
plot v(B0) v(B1)+2 v(B2)+4 v(B3)+6
* plot v(A0B0) v(A1B1)+2 v(A2B2)+4 v(A3B3)+6
plot v(A_IS_EQUAL_B)
* plot v(A3_B3NOT) v(A2_B2NOT_A3B3XNOR)+2 v(A1_B1NOT_A3B3XNOR_A2B2XOR)+4 v(A0_B0NOT_A3B3XNOR_A2B2XOR_A1B1XOR)+6
plot v(A_greater_than_B)
* plot v(A3NOT_B3) v(A2NOT_B2_A3B3XNOR)+2 v(A1NOTB1_A2XNORB2_A3XNORB3)+4 v(A0NOTB0_A1XNORB1_A2XNORB2_A3XNORB3)+6
plot v(A_less_than_B)
* hardcopy image.ps v(node_a) v(node_b)+2 v(OUT)+4
.end
.endc