.include TSMC_180nm.txt
.include NAND.sub
.include NOT.sub
.include AND.sub
.include OR.sub
.include XOR.sub


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 node_a0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)

V_in_b0 node_b0 gnd PULSE(0 1.8 50ns 100ps 100ps 50ns 100ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 100ns 100ps 100ps 100ns 200ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 200ns 100ps 100ps 200ns 400ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 400ns 100ps 100ps 500ns 1000ns)

* V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
* V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 140ns)
* V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
* V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)


X1 node_a node_b node_c node_x gnd XOR
X2 node_c node_c_in node_sum node_x gnd XOR
X3 node_a node_b node_d node_x gnd AND
X4 node_c node_c_in node_e node_x gnd AND
X5 node_d node_e node_cout node_x gnd OR
C1 node_out gnd 100f


.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
* plot v(node_a) v(node_b)+2 v(node_out)+4 v(node_out_final)+6
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4 v(node_out_final)+6
plot v(node_a) v(node_b)+2 v(node_c_in)+4 v(node_sum)+6 v(node_cout)+8
hardcopy image.ps v(node_a) v(node_b)+2 v(node_c_in)+4 v(node_sum)+6 v(node_cout)+8
.end
.endc